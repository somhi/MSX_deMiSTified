library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f0f6c287",
    12 => x"86c0c64e",
    13 => x"49f0f6c2",
    14 => x"48d0e2c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087eee1",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48111e4f",
    50 => x"7808d4ff",
    51 => x"c14866c4",
    52 => x"58a6c888",
    53 => x"ed059870",
    54 => x"1e4f2687",
    55 => x"c348d4ff",
    56 => x"516878ff",
    57 => x"c14866c4",
    58 => x"58a6c888",
    59 => x"eb059870",
    60 => x"1e4f2687",
    61 => x"d4ff1e73",
    62 => x"7bffc34b",
    63 => x"ffc34a6b",
    64 => x"c8496b7b",
    65 => x"c3b17232",
    66 => x"4a6b7bff",
    67 => x"b27131c8",
    68 => x"6b7bffc3",
    69 => x"7232c849",
    70 => x"c44871b1",
    71 => x"264d2687",
    72 => x"264b264c",
    73 => x"5b5e0e4f",
    74 => x"710e5d5c",
    75 => x"4cd4ff4a",
    76 => x"ffc34972",
    77 => x"c27c7199",
    78 => x"05bfd0e2",
    79 => x"66d087c8",
    80 => x"d430c948",
    81 => x"66d058a6",
    82 => x"c329d849",
    83 => x"7c7199ff",
    84 => x"d04966d0",
    85 => x"99ffc329",
    86 => x"66d07c71",
    87 => x"c329c849",
    88 => x"7c7199ff",
    89 => x"c34966d0",
    90 => x"7c7199ff",
    91 => x"29d04972",
    92 => x"7199ffc3",
    93 => x"c94b6c7c",
    94 => x"c34dfff0",
    95 => x"d005abff",
    96 => x"7cffc387",
    97 => x"8dc14b6c",
    98 => x"c387c602",
    99 => x"f002abff",
   100 => x"fe487387",
   101 => x"c01e87c7",
   102 => x"48d4ff49",
   103 => x"c178ffc3",
   104 => x"b7c8c381",
   105 => x"87f104a9",
   106 => x"731e4f26",
   107 => x"c487e71e",
   108 => x"c04bdff8",
   109 => x"f0ffc01e",
   110 => x"fd49f7c1",
   111 => x"86c487e7",
   112 => x"c005a8c1",
   113 => x"d4ff87ea",
   114 => x"78ffc348",
   115 => x"c0c0c0c1",
   116 => x"c01ec0c0",
   117 => x"e9c1f0e1",
   118 => x"87c9fd49",
   119 => x"987086c4",
   120 => x"ff87ca05",
   121 => x"ffc348d4",
   122 => x"cb48c178",
   123 => x"87e6fe87",
   124 => x"fe058bc1",
   125 => x"48c087fd",
   126 => x"1e87e6fc",
   127 => x"d4ff1e73",
   128 => x"78ffc348",
   129 => x"1ec04bd3",
   130 => x"c1f0ffc0",
   131 => x"d4fc49c1",
   132 => x"7086c487",
   133 => x"87ca0598",
   134 => x"c348d4ff",
   135 => x"48c178ff",
   136 => x"f1fd87cb",
   137 => x"058bc187",
   138 => x"c087dbff",
   139 => x"87f1fb48",
   140 => x"5c5b5e0e",
   141 => x"4cd4ff0e",
   142 => x"c687dbfd",
   143 => x"e1c01eea",
   144 => x"49c8c1f0",
   145 => x"c487defb",
   146 => x"02a8c186",
   147 => x"eafe87c8",
   148 => x"c148c087",
   149 => x"dafa87e2",
   150 => x"cf497087",
   151 => x"c699ffff",
   152 => x"c802a9ea",
   153 => x"87d3fe87",
   154 => x"cbc148c0",
   155 => x"7cffc387",
   156 => x"fc4bf1c0",
   157 => x"987087f4",
   158 => x"87ebc002",
   159 => x"ffc01ec0",
   160 => x"49fac1f0",
   161 => x"c487defa",
   162 => x"05987086",
   163 => x"ffc387d9",
   164 => x"c3496c7c",
   165 => x"7c7c7cff",
   166 => x"99c0c17c",
   167 => x"c187c402",
   168 => x"c087d548",
   169 => x"c287d148",
   170 => x"87c405ab",
   171 => x"87c848c0",
   172 => x"fe058bc1",
   173 => x"48c087fd",
   174 => x"1e87e4f9",
   175 => x"e2c21e73",
   176 => x"78c148d0",
   177 => x"d0ff4bc7",
   178 => x"fb78c248",
   179 => x"d0ff87c8",
   180 => x"c078c348",
   181 => x"d0e5c01e",
   182 => x"f949c0c1",
   183 => x"86c487c7",
   184 => x"c105a8c1",
   185 => x"abc24b87",
   186 => x"c087c505",
   187 => x"87f9c048",
   188 => x"ff058bc1",
   189 => x"f7fc87d0",
   190 => x"d4e2c287",
   191 => x"05987058",
   192 => x"1ec187cd",
   193 => x"c1f0ffc0",
   194 => x"d8f849d0",
   195 => x"ff86c487",
   196 => x"ffc348d4",
   197 => x"87e0c478",
   198 => x"58d8e2c2",
   199 => x"c248d0ff",
   200 => x"48d4ff78",
   201 => x"c178ffc3",
   202 => x"87f5f748",
   203 => x"5c5b5e0e",
   204 => x"4a710e5d",
   205 => x"ff4dffc3",
   206 => x"7c754cd4",
   207 => x"c448d0ff",
   208 => x"7c7578c3",
   209 => x"ffc01e72",
   210 => x"49d8c1f0",
   211 => x"c487d6f7",
   212 => x"02987086",
   213 => x"48c087c5",
   214 => x"7587f0c0",
   215 => x"7cfec37c",
   216 => x"d41ec0c8",
   217 => x"dcf54966",
   218 => x"7586c487",
   219 => x"757c757c",
   220 => x"e0dad87c",
   221 => x"6c7c754b",
   222 => x"c5059949",
   223 => x"058bc187",
   224 => x"7c7587f3",
   225 => x"c248d0ff",
   226 => x"f648c178",
   227 => x"ff1e87cf",
   228 => x"d0ff4ad4",
   229 => x"78d1c448",
   230 => x"c17affc3",
   231 => x"87f80589",
   232 => x"731e4f26",
   233 => x"c54b711e",
   234 => x"4adfcdee",
   235 => x"c348d4ff",
   236 => x"486878ff",
   237 => x"02a8fec3",
   238 => x"8ac187c5",
   239 => x"7287ed05",
   240 => x"87c5059a",
   241 => x"eac048c0",
   242 => x"029b7387",
   243 => x"66c887cc",
   244 => x"f449731e",
   245 => x"86c487c5",
   246 => x"66c887c6",
   247 => x"87eefe49",
   248 => x"c348d4ff",
   249 => x"737878ff",
   250 => x"87c5059b",
   251 => x"d048d0ff",
   252 => x"f448c178",
   253 => x"731e87eb",
   254 => x"c04a711e",
   255 => x"48d4ff4b",
   256 => x"ff78ffc3",
   257 => x"c3c448d0",
   258 => x"48d4ff78",
   259 => x"7278ffc3",
   260 => x"f0ffc01e",
   261 => x"f449d1c1",
   262 => x"86c487cb",
   263 => x"cd059870",
   264 => x"1ec0c887",
   265 => x"fd4966cc",
   266 => x"86c487f8",
   267 => x"d0ff4b70",
   268 => x"7378c248",
   269 => x"87e9f348",
   270 => x"5c5b5e0e",
   271 => x"1ec00e5d",
   272 => x"c1f0ffc0",
   273 => x"dcf349c9",
   274 => x"c21ed287",
   275 => x"fd49d8e2",
   276 => x"86c887d0",
   277 => x"84c14cc0",
   278 => x"04acb7d2",
   279 => x"e2c287f8",
   280 => x"49bf97d8",
   281 => x"c199c0c3",
   282 => x"c005a9c0",
   283 => x"e2c287e7",
   284 => x"49bf97df",
   285 => x"e2c231d0",
   286 => x"4abf97e0",
   287 => x"b17232c8",
   288 => x"97e1e2c2",
   289 => x"71b14abf",
   290 => x"ffffcf4c",
   291 => x"84c19cff",
   292 => x"e7c134ca",
   293 => x"e1e2c287",
   294 => x"c149bf97",
   295 => x"c299c631",
   296 => x"bf97e2e2",
   297 => x"2ab7c74a",
   298 => x"e2c2b172",
   299 => x"4abf97dd",
   300 => x"c29dcf4d",
   301 => x"bf97dee2",
   302 => x"ca9ac34a",
   303 => x"dfe2c232",
   304 => x"c24bbf97",
   305 => x"c2b27333",
   306 => x"bf97e0e2",
   307 => x"9bc0c34b",
   308 => x"732bb7c6",
   309 => x"c181c2b2",
   310 => x"70307148",
   311 => x"7548c149",
   312 => x"724d7030",
   313 => x"7184c14c",
   314 => x"b7c0c894",
   315 => x"87cc06ad",
   316 => x"2db734c1",
   317 => x"adb7c0c8",
   318 => x"87f4ff01",
   319 => x"dcf04874",
   320 => x"5b5e0e87",
   321 => x"f80e5d5c",
   322 => x"feeac286",
   323 => x"c278c048",
   324 => x"c01ef6e2",
   325 => x"87defb49",
   326 => x"987086c4",
   327 => x"c087c505",
   328 => x"87cec948",
   329 => x"7ec14dc0",
   330 => x"bfd0f8c0",
   331 => x"ece3c249",
   332 => x"4bc8714a",
   333 => x"7087f3ec",
   334 => x"87c20598",
   335 => x"f8c07ec0",
   336 => x"c249bfcc",
   337 => x"714ac8e4",
   338 => x"ddec4bc8",
   339 => x"05987087",
   340 => x"7ec087c2",
   341 => x"fdc0026e",
   342 => x"fce9c287",
   343 => x"eac24dbf",
   344 => x"7ebf9ff4",
   345 => x"ead6c548",
   346 => x"87c705a8",
   347 => x"bffce9c2",
   348 => x"6e87ce4d",
   349 => x"d5e9ca48",
   350 => x"87c502a8",
   351 => x"f1c748c0",
   352 => x"f6e2c287",
   353 => x"f949751e",
   354 => x"86c487ec",
   355 => x"c5059870",
   356 => x"c748c087",
   357 => x"f8c087dc",
   358 => x"c249bfcc",
   359 => x"714ac8e4",
   360 => x"c5eb4bc8",
   361 => x"05987087",
   362 => x"eac287c8",
   363 => x"78c148fe",
   364 => x"f8c087da",
   365 => x"c249bfd0",
   366 => x"714aece3",
   367 => x"e9ea4bc8",
   368 => x"02987087",
   369 => x"c087c5c0",
   370 => x"87e6c648",
   371 => x"97f4eac2",
   372 => x"d5c149bf",
   373 => x"cdc005a9",
   374 => x"f5eac287",
   375 => x"c249bf97",
   376 => x"c002a9ea",
   377 => x"48c087c5",
   378 => x"c287c7c6",
   379 => x"bf97f6e2",
   380 => x"e9c3487e",
   381 => x"cec002a8",
   382 => x"c3486e87",
   383 => x"c002a8eb",
   384 => x"48c087c5",
   385 => x"c287ebc5",
   386 => x"bf97c1e3",
   387 => x"c0059949",
   388 => x"e3c287cc",
   389 => x"49bf97c2",
   390 => x"c002a9c2",
   391 => x"48c087c5",
   392 => x"c287cfc5",
   393 => x"bf97c3e3",
   394 => x"faeac248",
   395 => x"484c7058",
   396 => x"eac288c1",
   397 => x"e3c258fe",
   398 => x"49bf97c4",
   399 => x"e3c28175",
   400 => x"4abf97c5",
   401 => x"a17232c8",
   402 => x"cbefc27e",
   403 => x"c2786e48",
   404 => x"bf97c6e3",
   405 => x"58a6c848",
   406 => x"bffeeac2",
   407 => x"87d4c202",
   408 => x"bfccf8c0",
   409 => x"c8e4c249",
   410 => x"4bc8714a",
   411 => x"7087fbe7",
   412 => x"c5c00298",
   413 => x"c348c087",
   414 => x"eac287f8",
   415 => x"c24cbff6",
   416 => x"c25cdfef",
   417 => x"bf97dbe3",
   418 => x"c231c849",
   419 => x"bf97dae3",
   420 => x"c249a14a",
   421 => x"bf97dce3",
   422 => x"7232d04a",
   423 => x"e3c249a1",
   424 => x"4abf97dd",
   425 => x"a17232d8",
   426 => x"9166c449",
   427 => x"bfcbefc2",
   428 => x"d3efc281",
   429 => x"e3e3c259",
   430 => x"c84abf97",
   431 => x"e2e3c232",
   432 => x"a24bbf97",
   433 => x"e4e3c24a",
   434 => x"d04bbf97",
   435 => x"4aa27333",
   436 => x"97e5e3c2",
   437 => x"9bcf4bbf",
   438 => x"a27333d8",
   439 => x"d7efc24a",
   440 => x"d3efc25a",
   441 => x"8ac24abf",
   442 => x"efc29274",
   443 => x"a17248d7",
   444 => x"87cac178",
   445 => x"97c8e3c2",
   446 => x"31c849bf",
   447 => x"97c7e3c2",
   448 => x"49a14abf",
   449 => x"59c6ebc2",
   450 => x"bfc2ebc2",
   451 => x"c731c549",
   452 => x"29c981ff",
   453 => x"59dfefc2",
   454 => x"97cde3c2",
   455 => x"32c84abf",
   456 => x"97cce3c2",
   457 => x"4aa24bbf",
   458 => x"6e9266c4",
   459 => x"dbefc282",
   460 => x"d3efc25a",
   461 => x"c278c048",
   462 => x"7248cfef",
   463 => x"efc278a1",
   464 => x"efc248df",
   465 => x"c278bfd3",
   466 => x"c248e3ef",
   467 => x"78bfd7ef",
   468 => x"bffeeac2",
   469 => x"87c9c002",
   470 => x"30c44874",
   471 => x"c9c07e70",
   472 => x"dbefc287",
   473 => x"30c448bf",
   474 => x"ebc27e70",
   475 => x"786e48c2",
   476 => x"8ef848c1",
   477 => x"4c264d26",
   478 => x"4f264b26",
   479 => x"5c5b5e0e",
   480 => x"4a710e5d",
   481 => x"bffeeac2",
   482 => x"7287cb02",
   483 => x"722bc74b",
   484 => x"9cffc14c",
   485 => x"4b7287c9",
   486 => x"4c722bc8",
   487 => x"c29cffc3",
   488 => x"83bfcbef",
   489 => x"bfc8f8c0",
   490 => x"87d902ab",
   491 => x"5bccf8c0",
   492 => x"1ef6e2c2",
   493 => x"fdf04973",
   494 => x"7086c487",
   495 => x"87c50598",
   496 => x"e6c048c0",
   497 => x"feeac287",
   498 => x"87d202bf",
   499 => x"91c44974",
   500 => x"81f6e2c2",
   501 => x"ffcf4d69",
   502 => x"9dffffff",
   503 => x"497487cb",
   504 => x"e2c291c2",
   505 => x"699f81f6",
   506 => x"fe48754d",
   507 => x"5e0e87c6",
   508 => x"0e5d5c5b",
   509 => x"c04d711e",
   510 => x"d049c11e",
   511 => x"86c487f2",
   512 => x"029c4c70",
   513 => x"c287c0c1",
   514 => x"754ac6eb",
   515 => x"87ffe049",
   516 => x"c0029870",
   517 => x"4a7487f1",
   518 => x"4bcb4975",
   519 => x"7087e5e1",
   520 => x"e2c00298",
   521 => x"741ec087",
   522 => x"87c7029c",
   523 => x"c048a6c4",
   524 => x"c487c578",
   525 => x"78c148a6",
   526 => x"cf4966c4",
   527 => x"86c487f2",
   528 => x"059c4c70",
   529 => x"7487c0ff",
   530 => x"e7fc2648",
   531 => x"5b5e0e87",
   532 => x"f80e5d5c",
   533 => x"9b4b7186",
   534 => x"c087c505",
   535 => x"87d4c248",
   536 => x"c04da3c8",
   537 => x"0266d87d",
   538 => x"66d887c7",
   539 => x"c505bf97",
   540 => x"c148c087",
   541 => x"66d887fe",
   542 => x"87f2fd49",
   543 => x"026e7e70",
   544 => x"6e87efc1",
   545 => x"6981dc49",
   546 => x"da496e7d",
   547 => x"4ca3c481",
   548 => x"c27c699f",
   549 => x"02bffeea",
   550 => x"496e87d0",
   551 => x"699f81d4",
   552 => x"ffc04a49",
   553 => x"32d09aff",
   554 => x"4ac087c2",
   555 => x"6c484972",
   556 => x"c07c7080",
   557 => x"49a3cc7b",
   558 => x"a3d0796c",
   559 => x"c479c049",
   560 => x"78c048a6",
   561 => x"c44aa3d4",
   562 => x"91c84966",
   563 => x"c049a172",
   564 => x"c4796c41",
   565 => x"80c14866",
   566 => x"c458a6c8",
   567 => x"ff04a8b7",
   568 => x"4a6d87e2",
   569 => x"2ac52ac9",
   570 => x"49a3f4c0",
   571 => x"486e7972",
   572 => x"48c087c2",
   573 => x"fbf98ef8",
   574 => x"5b5e0e87",
   575 => x"710e5d5c",
   576 => x"c8f8c04c",
   577 => x"7478ff48",
   578 => x"cac1029c",
   579 => x"49a4c887",
   580 => x"c2c10269",
   581 => x"4a66d087",
   582 => x"d482496c",
   583 => x"66d05aa6",
   584 => x"eac2b94d",
   585 => x"ff4abffa",
   586 => x"719972ba",
   587 => x"e4c00299",
   588 => x"4ba4c487",
   589 => x"c3f9496b",
   590 => x"c27b7087",
   591 => x"49bff6ea",
   592 => x"7c71816c",
   593 => x"eac2b975",
   594 => x"ff4abffa",
   595 => x"719972ba",
   596 => x"dcff0599",
   597 => x"f87c7587",
   598 => x"731e87da",
   599 => x"9b4b711e",
   600 => x"c887c702",
   601 => x"056949a3",
   602 => x"48c087c5",
   603 => x"c287ebc0",
   604 => x"4abfcfef",
   605 => x"6949a3c4",
   606 => x"c289c249",
   607 => x"91bff6ea",
   608 => x"c24aa271",
   609 => x"49bffaea",
   610 => x"a271996b",
   611 => x"1e66c84a",
   612 => x"e1e94972",
   613 => x"7086c487",
   614 => x"dbf74849",
   615 => x"1e731e87",
   616 => x"029b4b71",
   617 => x"a3c887c7",
   618 => x"c5056949",
   619 => x"c048c087",
   620 => x"efc287eb",
   621 => x"c44abfcf",
   622 => x"496949a3",
   623 => x"eac289c2",
   624 => x"7191bff6",
   625 => x"eac24aa2",
   626 => x"6b49bffa",
   627 => x"4aa27199",
   628 => x"721e66c8",
   629 => x"87d4e549",
   630 => x"497086c4",
   631 => x"87d8f648",
   632 => x"5c5b5e0e",
   633 => x"86f80e5d",
   634 => x"a6c44b71",
   635 => x"c878ff48",
   636 => x"4d6949a3",
   637 => x"a3d44cc0",
   638 => x"c849744a",
   639 => x"49a17291",
   640 => x"66d84969",
   641 => x"70887148",
   642 => x"a966d87e",
   643 => x"6e87ca01",
   644 => x"87c506ad",
   645 => x"6e5ca6c8",
   646 => x"c484c14d",
   647 => x"ff04acb7",
   648 => x"486687d4",
   649 => x"cbf58ef8",
   650 => x"5b5e0e87",
   651 => x"ec0e5d5c",
   652 => x"59a6c886",
   653 => x"c148a6c8",
   654 => x"ffffffff",
   655 => x"80c478ff",
   656 => x"4dc078ff",
   657 => x"66c44cc0",
   658 => x"7483d44b",
   659 => x"7391c849",
   660 => x"4a7549a1",
   661 => x"a27392c8",
   662 => x"6e49697e",
   663 => x"a6d489bf",
   664 => x"05ad7459",
   665 => x"a6d087c6",
   666 => x"78bf6e48",
   667 => x"c04866d0",
   668 => x"cf04a8b7",
   669 => x"4966d087",
   670 => x"03a966c8",
   671 => x"a6d087c6",
   672 => x"59a6cc5c",
   673 => x"b7c484c1",
   674 => x"f9fe04ac",
   675 => x"c485c187",
   676 => x"fe04adb7",
   677 => x"66cc87ee",
   678 => x"f38eec48",
   679 => x"5e0e87d6",
   680 => x"0e5d5c5b",
   681 => x"4b7186f0",
   682 => x"4c66e0c0",
   683 => x"9b732cc9",
   684 => x"87e1c302",
   685 => x"6949a3c8",
   686 => x"87d9c302",
   687 => x"c049a3d0",
   688 => x"6b7966e0",
   689 => x"c302ac7e",
   690 => x"eac287cb",
   691 => x"ff49bffa",
   692 => x"744a71b9",
   693 => x"6e48719a",
   694 => x"58a6cc98",
   695 => x"c44da3c4",
   696 => x"786d48a6",
   697 => x"05aa66c8",
   698 => x"7b7487c5",
   699 => x"7287d1c2",
   700 => x"fb49731e",
   701 => x"86c487ea",
   702 => x"c0487e70",
   703 => x"d004a8b7",
   704 => x"4aa3d487",
   705 => x"91c8496e",
   706 => x"2149a172",
   707 => x"c77d697b",
   708 => x"cc7bc087",
   709 => x"7d6949a3",
   710 => x"731e66c8",
   711 => x"87c0fb49",
   712 => x"7e7086c4",
   713 => x"49a3f4c0",
   714 => x"6948a6cc",
   715 => x"4866c878",
   716 => x"06a866cc",
   717 => x"486e87c9",
   718 => x"04a8b7c0",
   719 => x"6e87e0c0",
   720 => x"a8b7c048",
   721 => x"87ecc004",
   722 => x"6e4aa3d4",
   723 => x"7291c849",
   724 => x"66c849a1",
   725 => x"70886948",
   726 => x"a966cc49",
   727 => x"7387d506",
   728 => x"87c5fb49",
   729 => x"a3d44970",
   730 => x"7291c84a",
   731 => x"66c849a1",
   732 => x"7966c441",
   733 => x"49748c6b",
   734 => x"f549731e",
   735 => x"86c487fb",
   736 => x"4966e0c0",
   737 => x"0299ffc7",
   738 => x"e2c287cb",
   739 => x"49731ef6",
   740 => x"c487c7f7",
   741 => x"ef8ef086",
   742 => x"731e87da",
   743 => x"9b4b711e",
   744 => x"87e4c002",
   745 => x"5be3efc2",
   746 => x"8ac24a73",
   747 => x"bff6eac2",
   748 => x"efc29249",
   749 => x"7248bfcf",
   750 => x"e7efc280",
   751 => x"c4487158",
   752 => x"c6ebc230",
   753 => x"87edc058",
   754 => x"48dfefc2",
   755 => x"bfd3efc2",
   756 => x"e3efc278",
   757 => x"d7efc248",
   758 => x"eac278bf",
   759 => x"c902bffe",
   760 => x"f6eac287",
   761 => x"31c449bf",
   762 => x"efc287c7",
   763 => x"c449bfdb",
   764 => x"c6ebc231",
   765 => x"87c0ee59",
   766 => x"5c5b5e0e",
   767 => x"c04a710e",
   768 => x"029a724b",
   769 => x"da87e1c0",
   770 => x"699f49a2",
   771 => x"feeac24b",
   772 => x"87cf02bf",
   773 => x"9f49a2d4",
   774 => x"c04c4969",
   775 => x"d09cffff",
   776 => x"c087c234",
   777 => x"b349744c",
   778 => x"edfd4973",
   779 => x"87c6ed87",
   780 => x"5c5b5e0e",
   781 => x"86f40e5d",
   782 => x"7ec04a71",
   783 => x"d8029a72",
   784 => x"f2e2c287",
   785 => x"c278c048",
   786 => x"c248eae2",
   787 => x"78bfe3ef",
   788 => x"48eee2c2",
   789 => x"bfdfefc2",
   790 => x"d3ebc278",
   791 => x"c250c048",
   792 => x"49bfc2eb",
   793 => x"bff2e2c2",
   794 => x"03aa714a",
   795 => x"7287c0c4",
   796 => x"0599cf49",
   797 => x"c287e1c0",
   798 => x"c21ef6e2",
   799 => x"49bfeae2",
   800 => x"48eae2c2",
   801 => x"7178a1c1",
   802 => x"87eaddff",
   803 => x"f8c086c4",
   804 => x"e2c248c4",
   805 => x"87cc78f6",
   806 => x"bfc4f8c0",
   807 => x"80e0c048",
   808 => x"58c8f8c0",
   809 => x"bff2e2c2",
   810 => x"c280c148",
   811 => x"2758f6e2",
   812 => x"00000e04",
   813 => x"4dbf97bf",
   814 => x"e2c2029d",
   815 => x"ade5c387",
   816 => x"87dbc202",
   817 => x"bfc4f8c0",
   818 => x"49a3cb4b",
   819 => x"accf4c11",
   820 => x"87d2c105",
   821 => x"99df4975",
   822 => x"91cd89c1",
   823 => x"81c6ebc2",
   824 => x"124aa3c1",
   825 => x"4aa3c351",
   826 => x"a3c55112",
   827 => x"c751124a",
   828 => x"51124aa3",
   829 => x"124aa3c9",
   830 => x"4aa3ce51",
   831 => x"a3d05112",
   832 => x"d251124a",
   833 => x"51124aa3",
   834 => x"124aa3d4",
   835 => x"4aa3d651",
   836 => x"a3d85112",
   837 => x"dc51124a",
   838 => x"51124aa3",
   839 => x"124aa3de",
   840 => x"c07ec151",
   841 => x"497487f9",
   842 => x"c00599c8",
   843 => x"497487ea",
   844 => x"d00599d0",
   845 => x"0266dc87",
   846 => x"7387cac0",
   847 => x"0f66dc49",
   848 => x"d3029870",
   849 => x"c0056e87",
   850 => x"ebc287c6",
   851 => x"50c048c6",
   852 => x"bfc4f8c0",
   853 => x"87e7c248",
   854 => x"48d3ebc2",
   855 => x"c27e50c0",
   856 => x"49bfc2eb",
   857 => x"bff2e2c2",
   858 => x"04aa714a",
   859 => x"c287c0fc",
   860 => x"05bfe3ef",
   861 => x"c287c8c0",
   862 => x"02bffeea",
   863 => x"c087fec1",
   864 => x"ff48c8f8",
   865 => x"eee2c278",
   866 => x"efe749bf",
   867 => x"c2497087",
   868 => x"c459f2e2",
   869 => x"e2c248a6",
   870 => x"c278bfee",
   871 => x"02bffeea",
   872 => x"c487d8c0",
   873 => x"ffcf4966",
   874 => x"99f8ffff",
   875 => x"c5c002a9",
   876 => x"c04dc087",
   877 => x"4dc187e1",
   878 => x"c487dcc0",
   879 => x"ffcf4966",
   880 => x"02a999f8",
   881 => x"c887c8c0",
   882 => x"78c048a6",
   883 => x"c887c5c0",
   884 => x"78c148a6",
   885 => x"754d66c8",
   886 => x"e0c0059d",
   887 => x"4966c487",
   888 => x"eac289c2",
   889 => x"914abff6",
   890 => x"bfcfefc2",
   891 => x"eae2c24a",
   892 => x"78a17248",
   893 => x"48f2e2c2",
   894 => x"e2f978c0",
   895 => x"f448c087",
   896 => x"87f0e58e",
   897 => x"00000000",
   898 => x"ffffffff",
   899 => x"00000e14",
   900 => x"00000e1d",
   901 => x"33544146",
   902 => x"20202032",
   903 => x"54414600",
   904 => x"20203631",
   905 => x"ff1e0020",
   906 => x"ffc348d4",
   907 => x"26486878",
   908 => x"d4ff1e4f",
   909 => x"78ffc348",
   910 => x"c848d0ff",
   911 => x"d4ff78e1",
   912 => x"c278d448",
   913 => x"ff48e7ef",
   914 => x"2650bfd4",
   915 => x"d0ff1e4f",
   916 => x"78e0c048",
   917 => x"ff1e4f26",
   918 => x"497087cc",
   919 => x"87c60299",
   920 => x"05a9fbc0",
   921 => x"487187f1",
   922 => x"5e0e4f26",
   923 => x"710e5c5b",
   924 => x"fe4cc04b",
   925 => x"497087f0",
   926 => x"f9c00299",
   927 => x"a9ecc087",
   928 => x"87f2c002",
   929 => x"02a9fbc0",
   930 => x"cc87ebc0",
   931 => x"03acb766",
   932 => x"66d087c7",
   933 => x"7187c202",
   934 => x"02997153",
   935 => x"84c187c2",
   936 => x"7087c3fe",
   937 => x"cd029949",
   938 => x"a9ecc087",
   939 => x"c087c702",
   940 => x"ff05a9fb",
   941 => x"66d087d5",
   942 => x"c087c302",
   943 => x"ecc07b97",
   944 => x"87c405a9",
   945 => x"87c54a74",
   946 => x"0ac04a74",
   947 => x"c248728a",
   948 => x"264d2687",
   949 => x"264b264c",
   950 => x"c9fd1e4f",
   951 => x"c0497087",
   952 => x"04a9b7f0",
   953 => x"f9c087ca",
   954 => x"c301a9b7",
   955 => x"89f0c087",
   956 => x"a9b7c1c1",
   957 => x"c187ca04",
   958 => x"01a9b7da",
   959 => x"f7c087c3",
   960 => x"26487189",
   961 => x"5b5e0e4f",
   962 => x"4a710e5c",
   963 => x"724cd4ff",
   964 => x"87eac049",
   965 => x"029b4b70",
   966 => x"8bc187c2",
   967 => x"c848d0ff",
   968 => x"d5c178c5",
   969 => x"c649737c",
   970 => x"fae0c231",
   971 => x"484abf97",
   972 => x"7c70b071",
   973 => x"c448d0ff",
   974 => x"fe487378",
   975 => x"5e0e87d5",
   976 => x"0e5d5c5b",
   977 => x"4c7186f8",
   978 => x"e4fb7ec0",
   979 => x"c04bc087",
   980 => x"bf97ebff",
   981 => x"04a9c049",
   982 => x"f9fb87cf",
   983 => x"c083c187",
   984 => x"bf97ebff",
   985 => x"f106ab49",
   986 => x"ebffc087",
   987 => x"cf02bf97",
   988 => x"87f2fa87",
   989 => x"02994970",
   990 => x"ecc087c6",
   991 => x"87f105a9",
   992 => x"e1fa4bc0",
   993 => x"fa4d7087",
   994 => x"a6c887dc",
   995 => x"87d6fa58",
   996 => x"83c14a70",
   997 => x"9749a4c8",
   998 => x"02ad4969",
   999 => x"ffc087c7",
  1000 => x"e7c005ad",
  1001 => x"49a4c987",
  1002 => x"c4496997",
  1003 => x"c702a966",
  1004 => x"ffc04887",
  1005 => x"87d405a8",
  1006 => x"9749a4ca",
  1007 => x"02aa4969",
  1008 => x"ffc087c6",
  1009 => x"87c405aa",
  1010 => x"87d07ec1",
  1011 => x"02adecc0",
  1012 => x"fbc087c6",
  1013 => x"87c405ad",
  1014 => x"7ec14bc0",
  1015 => x"e1fe026e",
  1016 => x"87e9f987",
  1017 => x"8ef84873",
  1018 => x"0087e6fb",
  1019 => x"5c5b5e0e",
  1020 => x"711e0e5d",
  1021 => x"4d4cc04b",
  1022 => x"e8c004ab",
  1023 => x"fefcc087",
  1024 => x"029d751e",
  1025 => x"4ac087c4",
  1026 => x"4ac187c2",
  1027 => x"dff04972",
  1028 => x"7086c487",
  1029 => x"6e84c17e",
  1030 => x"7387c205",
  1031 => x"7385c14c",
  1032 => x"d8ff06ac",
  1033 => x"26486e87",
  1034 => x"4c264d26",
  1035 => x"4f264b26",
  1036 => x"5c5b5e0e",
  1037 => x"711e0e5d",
  1038 => x"91de494c",
  1039 => x"4dc1f0c2",
  1040 => x"6d978571",
  1041 => x"87ddc102",
  1042 => x"bfecefc2",
  1043 => x"7282744a",
  1044 => x"87d8fe49",
  1045 => x"026e7e70",
  1046 => x"c287f3c0",
  1047 => x"6e4bf4ef",
  1048 => x"ff49cb4a",
  1049 => x"7487c1c1",
  1050 => x"c193cb4b",
  1051 => x"c483dde3",
  1052 => x"e9c2c183",
  1053 => x"c149747b",
  1054 => x"7587d1c3",
  1055 => x"c0f0c27b",
  1056 => x"1e49bf97",
  1057 => x"49f4efc2",
  1058 => x"87f0ddc1",
  1059 => x"497486c4",
  1060 => x"87f8c2c1",
  1061 => x"c4c149c0",
  1062 => x"efc287d7",
  1063 => x"78c048e8",
  1064 => x"cbdd49c1",
  1065 => x"fffd2687",
  1066 => x"616f4c87",
  1067 => x"676e6964",
  1068 => x"002e2e2e",
  1069 => x"5c5b5e0e",
  1070 => x"4a4b710e",
  1071 => x"bfecefc2",
  1072 => x"fc497282",
  1073 => x"4c7087e6",
  1074 => x"87c4029c",
  1075 => x"87e8ec49",
  1076 => x"48ecefc2",
  1077 => x"49c178c0",
  1078 => x"fd87d5dc",
  1079 => x"5e0e87cc",
  1080 => x"0e5d5c5b",
  1081 => x"e2c286f4",
  1082 => x"4cc04df6",
  1083 => x"c048a6c4",
  1084 => x"ecefc278",
  1085 => x"a9c049bf",
  1086 => x"87c1c106",
  1087 => x"48f6e2c2",
  1088 => x"f8c00298",
  1089 => x"fefcc087",
  1090 => x"0266c81e",
  1091 => x"a6c487c7",
  1092 => x"c578c048",
  1093 => x"48a6c487",
  1094 => x"66c478c1",
  1095 => x"87d0ec49",
  1096 => x"4d7086c4",
  1097 => x"66c484c1",
  1098 => x"c880c148",
  1099 => x"efc258a6",
  1100 => x"ac49bfec",
  1101 => x"7587c603",
  1102 => x"c8ff059d",
  1103 => x"754cc087",
  1104 => x"e0c3029d",
  1105 => x"fefcc087",
  1106 => x"0266c81e",
  1107 => x"a6cc87c7",
  1108 => x"c578c048",
  1109 => x"48a6cc87",
  1110 => x"66cc78c1",
  1111 => x"87d0eb49",
  1112 => x"7e7086c4",
  1113 => x"e9c2026e",
  1114 => x"cb496e87",
  1115 => x"49699781",
  1116 => x"c10299d0",
  1117 => x"c2c187d6",
  1118 => x"49744af4",
  1119 => x"e3c191cb",
  1120 => x"797281dd",
  1121 => x"ffc381c8",
  1122 => x"de497451",
  1123 => x"c1f0c291",
  1124 => x"c285714d",
  1125 => x"c17d97c1",
  1126 => x"e0c049a5",
  1127 => x"c6ebc251",
  1128 => x"d202bf97",
  1129 => x"c284c187",
  1130 => x"ebc24ba5",
  1131 => x"49db4ac6",
  1132 => x"87f4fbfe",
  1133 => x"cd87dbc1",
  1134 => x"51c049a5",
  1135 => x"a5c284c1",
  1136 => x"cb4a6e4b",
  1137 => x"dffbfe49",
  1138 => x"87c6c187",
  1139 => x"4af0c0c1",
  1140 => x"91cb4974",
  1141 => x"81dde3c1",
  1142 => x"ebc27972",
  1143 => x"02bf97c6",
  1144 => x"497487d8",
  1145 => x"84c191de",
  1146 => x"4bc1f0c2",
  1147 => x"ebc28371",
  1148 => x"49dd4ac6",
  1149 => x"87f0fafe",
  1150 => x"4b7487d8",
  1151 => x"f0c293de",
  1152 => x"a3cb83c1",
  1153 => x"c151c049",
  1154 => x"4a6e7384",
  1155 => x"fafe49cb",
  1156 => x"66c487d6",
  1157 => x"c880c148",
  1158 => x"acc758a6",
  1159 => x"87c5c003",
  1160 => x"e0fc056e",
  1161 => x"f4487487",
  1162 => x"87fcf78e",
  1163 => x"711e731e",
  1164 => x"91cb494b",
  1165 => x"81dde3c1",
  1166 => x"c24aa1c8",
  1167 => x"1248fae0",
  1168 => x"4aa1c950",
  1169 => x"48ebffc0",
  1170 => x"81ca5012",
  1171 => x"48c0f0c2",
  1172 => x"f0c25011",
  1173 => x"49bf97c0",
  1174 => x"c149c01e",
  1175 => x"c287ddd6",
  1176 => x"de48e8ef",
  1177 => x"d649c178",
  1178 => x"f62687c6",
  1179 => x"711e87fe",
  1180 => x"91cb494a",
  1181 => x"81dde3c1",
  1182 => x"481181c8",
  1183 => x"58ecefc2",
  1184 => x"48ecefc2",
  1185 => x"49c178c0",
  1186 => x"2687e5d5",
  1187 => x"49c01e4f",
  1188 => x"87ddfcc0",
  1189 => x"711e4f26",
  1190 => x"87d20299",
  1191 => x"48f2e4c1",
  1192 => x"80f750c0",
  1193 => x"40eec9c1",
  1194 => x"78d6e3c1",
  1195 => x"e4c187ce",
  1196 => x"e3c148ee",
  1197 => x"80fc78cf",
  1198 => x"78cdcac1",
  1199 => x"5e0e4f26",
  1200 => x"710e5c5b",
  1201 => x"92cb4a4c",
  1202 => x"82dde3c1",
  1203 => x"c949a2c8",
  1204 => x"6b974ba2",
  1205 => x"69971e4b",
  1206 => x"82ca1e49",
  1207 => x"e7c04912",
  1208 => x"49c087d8",
  1209 => x"7487c9d4",
  1210 => x"dff9c049",
  1211 => x"f48ef887",
  1212 => x"731e87f8",
  1213 => x"494b711e",
  1214 => x"7387c3ff",
  1215 => x"87fefe49",
  1216 => x"1e87e9f4",
  1217 => x"4b711e73",
  1218 => x"024aa3c6",
  1219 => x"8ac187db",
  1220 => x"8a87d602",
  1221 => x"87dac102",
  1222 => x"fcc0028a",
  1223 => x"c0028a87",
  1224 => x"028a87e1",
  1225 => x"dbc187cb",
  1226 => x"fd49c787",
  1227 => x"dec187c0",
  1228 => x"ecefc287",
  1229 => x"cbc102bf",
  1230 => x"88c14887",
  1231 => x"58f0efc2",
  1232 => x"c287c1c1",
  1233 => x"02bff0ef",
  1234 => x"c287f9c0",
  1235 => x"48bfecef",
  1236 => x"efc280c1",
  1237 => x"ebc058f0",
  1238 => x"ecefc287",
  1239 => x"89c649bf",
  1240 => x"59f0efc2",
  1241 => x"03a9b7c0",
  1242 => x"efc287da",
  1243 => x"78c048ec",
  1244 => x"efc287d2",
  1245 => x"cb02bff0",
  1246 => x"ecefc287",
  1247 => x"80c648bf",
  1248 => x"58f0efc2",
  1249 => x"e7d149c0",
  1250 => x"c0497387",
  1251 => x"f287fdf6",
  1252 => x"5e0e87da",
  1253 => x"710e5c5b",
  1254 => x"1e66cc4c",
  1255 => x"93cb4b74",
  1256 => x"83dde3c1",
  1257 => x"6a4aa3c4",
  1258 => x"cbf4fe49",
  1259 => x"ecc8c187",
  1260 => x"49a3c87b",
  1261 => x"c95166d4",
  1262 => x"66d849a3",
  1263 => x"49a3ca51",
  1264 => x"265166dc",
  1265 => x"0e87e3f1",
  1266 => x"5d5c5b5e",
  1267 => x"86d0ff0e",
  1268 => x"c459a6d8",
  1269 => x"78c048a6",
  1270 => x"c4c180c4",
  1271 => x"80c47866",
  1272 => x"80c478c1",
  1273 => x"efc278c1",
  1274 => x"78c148f0",
  1275 => x"bfe8efc2",
  1276 => x"05a8de48",
  1277 => x"e5f387cb",
  1278 => x"c8497087",
  1279 => x"f8ce59a6",
  1280 => x"87ede887",
  1281 => x"e887cfe9",
  1282 => x"4c7087dc",
  1283 => x"02acfbc0",
  1284 => x"d487d0c1",
  1285 => x"c2c10566",
  1286 => x"1e1ec087",
  1287 => x"e5c11ec1",
  1288 => x"49c01ed0",
  1289 => x"c187ebfd",
  1290 => x"c44a66d0",
  1291 => x"c7496a82",
  1292 => x"c1517481",
  1293 => x"6a1ed81e",
  1294 => x"e881c849",
  1295 => x"86d887ec",
  1296 => x"4866c4c1",
  1297 => x"c701a8c0",
  1298 => x"48a6c487",
  1299 => x"87ce78c1",
  1300 => x"4866c4c1",
  1301 => x"a6cc88c1",
  1302 => x"e787c358",
  1303 => x"a6cc87f8",
  1304 => x"7478c248",
  1305 => x"cccd029c",
  1306 => x"4866c487",
  1307 => x"a866c8c1",
  1308 => x"87c1cd03",
  1309 => x"c048a6d8",
  1310 => x"87eae678",
  1311 => x"d0c14c70",
  1312 => x"d6c205ac",
  1313 => x"7e66d887",
  1314 => x"7087cee9",
  1315 => x"59a6dc49",
  1316 => x"7087d3e6",
  1317 => x"acecc04c",
  1318 => x"87eac105",
  1319 => x"cb4966c4",
  1320 => x"66c0c191",
  1321 => x"4aa1c481",
  1322 => x"a1c84d6a",
  1323 => x"5266d84a",
  1324 => x"79eec9c1",
  1325 => x"7087efe5",
  1326 => x"d8029c4c",
  1327 => x"acfbc087",
  1328 => x"7487d202",
  1329 => x"87dee555",
  1330 => x"029c4c70",
  1331 => x"fbc087c7",
  1332 => x"eeff05ac",
  1333 => x"55e0c087",
  1334 => x"c055c1c2",
  1335 => x"66d47d97",
  1336 => x"05a96e49",
  1337 => x"66c487db",
  1338 => x"a866c848",
  1339 => x"c487ca04",
  1340 => x"80c14866",
  1341 => x"c858a6c8",
  1342 => x"4866c887",
  1343 => x"a6cc88c1",
  1344 => x"87e2e458",
  1345 => x"d0c14c70",
  1346 => x"87c805ac",
  1347 => x"c14866d0",
  1348 => x"58a6d480",
  1349 => x"02acd0c1",
  1350 => x"dc87eafd",
  1351 => x"66d448a6",
  1352 => x"4866d878",
  1353 => x"05a866dc",
  1354 => x"c087dcc9",
  1355 => x"c048a6e0",
  1356 => x"80c478f0",
  1357 => x"c47866cc",
  1358 => x"7e78c080",
  1359 => x"fbc04874",
  1360 => x"a6f0c088",
  1361 => x"02987058",
  1362 => x"4887d7c8",
  1363 => x"f0c088cb",
  1364 => x"987058a6",
  1365 => x"87e9c002",
  1366 => x"c088c948",
  1367 => x"7058a6f0",
  1368 => x"e1c30298",
  1369 => x"88c44887",
  1370 => x"58a6f0c0",
  1371 => x"d6029870",
  1372 => x"88c14887",
  1373 => x"58a6f0c0",
  1374 => x"c3029870",
  1375 => x"dbc787c8",
  1376 => x"a6e0c087",
  1377 => x"cc78c048",
  1378 => x"80c14866",
  1379 => x"e258a6d0",
  1380 => x"4c7087d4",
  1381 => x"02acecc0",
  1382 => x"e0c087d5",
  1383 => x"87c60266",
  1384 => x"5ca6e4c0",
  1385 => x"487487c9",
  1386 => x"c088f0c0",
  1387 => x"c058a6e8",
  1388 => x"cc02acec",
  1389 => x"87eee187",
  1390 => x"ecc04c70",
  1391 => x"f4ff05ac",
  1392 => x"66e0c087",
  1393 => x"4966d41e",
  1394 => x"66ecc01e",
  1395 => x"d0e5c11e",
  1396 => x"4966d41e",
  1397 => x"c087fbf6",
  1398 => x"dc1eca1e",
  1399 => x"91cb4966",
  1400 => x"8166d8c1",
  1401 => x"c448a6d8",
  1402 => x"66d878a1",
  1403 => x"f9e149bf",
  1404 => x"c086d887",
  1405 => x"c106a8b7",
  1406 => x"1ec187c7",
  1407 => x"66c81ede",
  1408 => x"e5e149bf",
  1409 => x"7086c887",
  1410 => x"08c04849",
  1411 => x"a6e4c088",
  1412 => x"a8b7c058",
  1413 => x"87e9c006",
  1414 => x"4866e0c0",
  1415 => x"03a8b7dd",
  1416 => x"bf6e87df",
  1417 => x"66e0c049",
  1418 => x"51e0c081",
  1419 => x"81c14966",
  1420 => x"c281bf6e",
  1421 => x"e0c051c1",
  1422 => x"81c24966",
  1423 => x"c081bf6e",
  1424 => x"c47ec151",
  1425 => x"d0e287dc",
  1426 => x"a6e4c087",
  1427 => x"87c9e258",
  1428 => x"58a6e8c0",
  1429 => x"05a8ecc0",
  1430 => x"c087cbc0",
  1431 => x"c048a6e4",
  1432 => x"c07866e0",
  1433 => x"deff87c4",
  1434 => x"66c487fc",
  1435 => x"c191cb49",
  1436 => x"714866c0",
  1437 => x"6e7e7080",
  1438 => x"6e82c84a",
  1439 => x"c081ca49",
  1440 => x"c05166e0",
  1441 => x"c14966e4",
  1442 => x"66e0c081",
  1443 => x"7148c189",
  1444 => x"c1497030",
  1445 => x"7a977189",
  1446 => x"bfddf3c2",
  1447 => x"66e0c049",
  1448 => x"4a6a9729",
  1449 => x"c0987148",
  1450 => x"6e58a6f0",
  1451 => x"6981c449",
  1452 => x"4866dc4d",
  1453 => x"02a866d8",
  1454 => x"d887c8c0",
  1455 => x"78c048a6",
  1456 => x"d887c5c0",
  1457 => x"78c148a6",
  1458 => x"c01e66d8",
  1459 => x"49751ee0",
  1460 => x"87d6deff",
  1461 => x"4c7086c8",
  1462 => x"06acb7c0",
  1463 => x"7487d4c1",
  1464 => x"49e0c085",
  1465 => x"4b758974",
  1466 => x"4aeddfc1",
  1467 => x"f7e6fe71",
  1468 => x"c085c287",
  1469 => x"c14866e8",
  1470 => x"a6ecc080",
  1471 => x"66ecc058",
  1472 => x"7081c149",
  1473 => x"c8c002a9",
  1474 => x"48a6d887",
  1475 => x"c5c078c0",
  1476 => x"48a6d887",
  1477 => x"66d878c1",
  1478 => x"49a4c21e",
  1479 => x"7148e0c0",
  1480 => x"1e497088",
  1481 => x"ddff4975",
  1482 => x"86c887c0",
  1483 => x"01a8b7c0",
  1484 => x"c087c0ff",
  1485 => x"c00266e8",
  1486 => x"496e87d1",
  1487 => x"e8c081c9",
  1488 => x"486e5166",
  1489 => x"78fecac1",
  1490 => x"6e87ccc0",
  1491 => x"c281c949",
  1492 => x"c1486e51",
  1493 => x"c178f2cb",
  1494 => x"87c6c07e",
  1495 => x"87f6dbff",
  1496 => x"026e4c70",
  1497 => x"c487f5c0",
  1498 => x"66c84866",
  1499 => x"cbc004a8",
  1500 => x"4866c487",
  1501 => x"a6c880c1",
  1502 => x"87e0c058",
  1503 => x"c14866c8",
  1504 => x"58a6cc88",
  1505 => x"c187d5c0",
  1506 => x"c005acc6",
  1507 => x"66cc87c8",
  1508 => x"d080c148",
  1509 => x"daff58a6",
  1510 => x"4c7087fc",
  1511 => x"c14866d0",
  1512 => x"58a6d480",
  1513 => x"c0029c74",
  1514 => x"66c487cb",
  1515 => x"66c8c148",
  1516 => x"fff204a8",
  1517 => x"d4daff87",
  1518 => x"4866c487",
  1519 => x"c003a8c7",
  1520 => x"efc287e5",
  1521 => x"78c048f0",
  1522 => x"cb4966c4",
  1523 => x"66c0c191",
  1524 => x"4aa1c481",
  1525 => x"52c04a6a",
  1526 => x"4866c479",
  1527 => x"a6c880c1",
  1528 => x"04a8c758",
  1529 => x"ff87dbff",
  1530 => x"fbe08ed0",
  1531 => x"00203a87",
  1532 => x"711e731e",
  1533 => x"c6029b4b",
  1534 => x"ecefc287",
  1535 => x"c778c048",
  1536 => x"ecefc21e",
  1537 => x"c11e49bf",
  1538 => x"c21edde3",
  1539 => x"49bfe8ef",
  1540 => x"cc87f4ee",
  1541 => x"e8efc286",
  1542 => x"f9e949bf",
  1543 => x"029b7387",
  1544 => x"e3c187c8",
  1545 => x"e5c049dd",
  1546 => x"dfff87f4",
  1547 => x"c21e87fe",
  1548 => x"c048fae0",
  1549 => x"c0e5c150",
  1550 => x"fbc049bf",
  1551 => x"48c087d1",
  1552 => x"c71e4f26",
  1553 => x"49c187e9",
  1554 => x"fe87e5fe",
  1555 => x"7087ece9",
  1556 => x"87cd0298",
  1557 => x"87e9f2fe",
  1558 => x"c4029870",
  1559 => x"c24ac187",
  1560 => x"724ac087",
  1561 => x"87ce059a",
  1562 => x"e2c11ec0",
  1563 => x"f0c049d6",
  1564 => x"86c487fb",
  1565 => x"ffc087fe",
  1566 => x"1ec087ea",
  1567 => x"49e1e2c1",
  1568 => x"87e9f0c0",
  1569 => x"e5fe1ec0",
  1570 => x"c0497087",
  1571 => x"c387def0",
  1572 => x"8ef887dc",
  1573 => x"44534f26",
  1574 => x"69616620",
  1575 => x"2e64656c",
  1576 => x"6f6f4200",
  1577 => x"676e6974",
  1578 => x"002e2e2e",
  1579 => x"c9e8c01e",
  1580 => x"eef3c087",
  1581 => x"2687f687",
  1582 => x"efc21e4f",
  1583 => x"78c048ec",
  1584 => x"48e8efc2",
  1585 => x"f9fd78c0",
  1586 => x"c087e187",
  1587 => x"804f2648",
  1588 => x"69784520",
  1589 => x"20800074",
  1590 => x"6b636142",
  1591 => x"00126e00",
  1592 => x"002c0100",
  1593 => x"00000000",
  1594 => x"0000126e",
  1595 => x"00002c1f",
  1596 => x"6e000000",
  1597 => x"3d000012",
  1598 => x"0000002c",
  1599 => x"126e0000",
  1600 => x"2c5b0000",
  1601 => x"00000000",
  1602 => x"00126e00",
  1603 => x"002c7900",
  1604 => x"00000000",
  1605 => x"0000126e",
  1606 => x"00002c97",
  1607 => x"6e000000",
  1608 => x"b5000012",
  1609 => x"0000002c",
  1610 => x"126e0000",
  1611 => x"00000000",
  1612 => x"00000000",
  1613 => x"00130300",
  1614 => x"00000000",
  1615 => x"00000000",
  1616 => x"00001944",
  1617 => x"544f4f42",
  1618 => x"20202020",
  1619 => x"004d4f52",
  1620 => x"64616f4c",
  1621 => x"002e2a20",
  1622 => x"48f0fe1e",
  1623 => x"09cd78c0",
  1624 => x"4f260979",
  1625 => x"f0fe1e1e",
  1626 => x"26487ebf",
  1627 => x"fe1e4f26",
  1628 => x"78c148f0",
  1629 => x"fe1e4f26",
  1630 => x"78c048f0",
  1631 => x"711e4f26",
  1632 => x"5252c04a",
  1633 => x"5e0e4f26",
  1634 => x"0e5d5c5b",
  1635 => x"4d7186f4",
  1636 => x"c17e6d97",
  1637 => x"6c974ca5",
  1638 => x"58a6c848",
  1639 => x"66c4486e",
  1640 => x"87c505a8",
  1641 => x"e6c048ff",
  1642 => x"87caff87",
  1643 => x"9749a5c2",
  1644 => x"a3714b6c",
  1645 => x"4b6b974b",
  1646 => x"6e7e6c97",
  1647 => x"c880c148",
  1648 => x"98c758a6",
  1649 => x"7058a6cc",
  1650 => x"e1fe7c97",
  1651 => x"f4487387",
  1652 => x"264d268e",
  1653 => x"264b264c",
  1654 => x"5b5e0e4f",
  1655 => x"86f40e5c",
  1656 => x"66d84c71",
  1657 => x"9affc34a",
  1658 => x"974ba4c2",
  1659 => x"a173496c",
  1660 => x"97517249",
  1661 => x"486e7e6c",
  1662 => x"a6c880c1",
  1663 => x"cc98c758",
  1664 => x"547058a6",
  1665 => x"caff8ef4",
  1666 => x"fd1e1e87",
  1667 => x"bfe087e8",
  1668 => x"e0c0494a",
  1669 => x"cb0299c0",
  1670 => x"c21e7287",
  1671 => x"fe49d3f3",
  1672 => x"86c487f7",
  1673 => x"7087fdfc",
  1674 => x"87c2fd7e",
  1675 => x"1e4f2626",
  1676 => x"49d3f3c2",
  1677 => x"c187c7fd",
  1678 => x"fc49c9e8",
  1679 => x"d9c587da",
  1680 => x"0e4f2687",
  1681 => x"5d5c5b5e",
  1682 => x"f2f3c20e",
  1683 => x"eac14abf",
  1684 => x"4c49bfd7",
  1685 => x"4d71bc72",
  1686 => x"c087dbfc",
  1687 => x"d049744b",
  1688 => x"87d50299",
  1689 => x"99d04975",
  1690 => x"1ec01e71",
  1691 => x"4ae9f0c1",
  1692 => x"49128273",
  1693 => x"c887e4c0",
  1694 => x"2d2cc186",
  1695 => x"04abc883",
  1696 => x"fb87daff",
  1697 => x"eac187e8",
  1698 => x"f3c248d7",
  1699 => x"2678bff2",
  1700 => x"264c264d",
  1701 => x"004f264b",
  1702 => x"1e000000",
  1703 => x"c848d0ff",
  1704 => x"d4ff78e1",
  1705 => x"c478c548",
  1706 => x"87c30266",
  1707 => x"c878e0c3",
  1708 => x"87c60266",
  1709 => x"c348d4ff",
  1710 => x"d4ff78f0",
  1711 => x"ff787148",
  1712 => x"e1c848d0",
  1713 => x"78e0c078",
  1714 => x"5e0e4f26",
  1715 => x"710e5c5b",
  1716 => x"d3f3c24c",
  1717 => x"87eefa49",
  1718 => x"b7c04a70",
  1719 => x"e3c204aa",
  1720 => x"aae0c387",
  1721 => x"c187c905",
  1722 => x"c148cdee",
  1723 => x"87d4c278",
  1724 => x"05aaf0c3",
  1725 => x"eec187c9",
  1726 => x"78c148c9",
  1727 => x"c187f5c1",
  1728 => x"02bfcdee",
  1729 => x"4b7287c7",
  1730 => x"c2b3c0c2",
  1731 => x"744b7287",
  1732 => x"87d1059c",
  1733 => x"bfc9eec1",
  1734 => x"cdeec11e",
  1735 => x"49721ebf",
  1736 => x"c887f8fd",
  1737 => x"c9eec186",
  1738 => x"e0c002bf",
  1739 => x"c4497387",
  1740 => x"c19129b7",
  1741 => x"7381e9ef",
  1742 => x"c29acf4a",
  1743 => x"7248c192",
  1744 => x"ff4a7030",
  1745 => x"694872ba",
  1746 => x"db797098",
  1747 => x"c4497387",
  1748 => x"c19129b7",
  1749 => x"7381e9ef",
  1750 => x"c29acf4a",
  1751 => x"7248c392",
  1752 => x"484a7030",
  1753 => x"7970b069",
  1754 => x"48cdeec1",
  1755 => x"eec178c0",
  1756 => x"78c048c9",
  1757 => x"49d3f3c2",
  1758 => x"7087cbf8",
  1759 => x"aab7c04a",
  1760 => x"87ddfd03",
  1761 => x"c8fc48c0",
  1762 => x"00000087",
  1763 => x"00000000",
  1764 => x"4a711e00",
  1765 => x"87f2fc49",
  1766 => x"c01e4f26",
  1767 => x"c449724a",
  1768 => x"e9efc191",
  1769 => x"c179c081",
  1770 => x"aab7d082",
  1771 => x"2687ee04",
  1772 => x"5b5e0e4f",
  1773 => x"710e5d5c",
  1774 => x"87faf64d",
  1775 => x"b7c44a75",
  1776 => x"efc1922a",
  1777 => x"4c7582e9",
  1778 => x"94c29ccf",
  1779 => x"744b496a",
  1780 => x"c29bc32b",
  1781 => x"70307448",
  1782 => x"74bcff4c",
  1783 => x"70987148",
  1784 => x"87caf67a",
  1785 => x"e6fa4873",
  1786 => x"00000087",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"00000000",
  1794 => x"00000000",
  1795 => x"00000000",
  1796 => x"00000000",
  1797 => x"00000000",
  1798 => x"00000000",
  1799 => x"00000000",
  1800 => x"00000000",
  1801 => x"00000000",
  1802 => x"261e1600",
  1803 => x"3d362e25",
  1804 => x"d0ff1e3e",
  1805 => x"78e1c848",
  1806 => x"d4ff4871",
  1807 => x"4f267808",
  1808 => x"48d0ff1e",
  1809 => x"7178e1c8",
  1810 => x"08d4ff48",
  1811 => x"4866c478",
  1812 => x"7808d4ff",
  1813 => x"711e4f26",
  1814 => x"4966c44a",
  1815 => x"ff49721e",
  1816 => x"d0ff87de",
  1817 => x"78e0c048",
  1818 => x"1e4f2626",
  1819 => x"66c44a71",
  1820 => x"a2e0c11e",
  1821 => x"87c8ff49",
  1822 => x"c84966c8",
  1823 => x"d4ff29b7",
  1824 => x"ff787148",
  1825 => x"e0c048d0",
  1826 => x"4f262678",
  1827 => x"4ad4ff1e",
  1828 => x"ff7affc3",
  1829 => x"e1c848d0",
  1830 => x"c27ade78",
  1831 => x"7abfddf3",
  1832 => x"28c84849",
  1833 => x"48717a70",
  1834 => x"7a7028d0",
  1835 => x"28d84871",
  1836 => x"d0ff7a70",
  1837 => x"78e0c048",
  1838 => x"5e0e4f26",
  1839 => x"0e5d5c5b",
  1840 => x"f3c24c71",
  1841 => x"4b4dbfdd",
  1842 => x"66d02b74",
  1843 => x"d483c19b",
  1844 => x"c204ab66",
  1845 => x"744bc087",
  1846 => x"4966d04a",
  1847 => x"b9ff3172",
  1848 => x"48739975",
  1849 => x"4a703072",
  1850 => x"c2b07148",
  1851 => x"fe58e1f3",
  1852 => x"4d2687da",
  1853 => x"4b264c26",
  1854 => x"ff1e4f26",
  1855 => x"c9c848d0",
  1856 => x"ff487178",
  1857 => x"267808d4",
  1858 => x"4a711e4f",
  1859 => x"ff87eb49",
  1860 => x"78c848d0",
  1861 => x"731e4f26",
  1862 => x"c24b711e",
  1863 => x"02bfedf3",
  1864 => x"ebc287c3",
  1865 => x"48d0ff87",
  1866 => x"7378c9c8",
  1867 => x"b1e0c049",
  1868 => x"7148d4ff",
  1869 => x"e1f3c278",
  1870 => x"c878c048",
  1871 => x"87c50266",
  1872 => x"c249ffc3",
  1873 => x"c249c087",
  1874 => x"cc59e9f3",
  1875 => x"87c60266",
  1876 => x"4ad5d5c5",
  1877 => x"ffcf87c4",
  1878 => x"f3c24aff",
  1879 => x"f3c25aed",
  1880 => x"78c148ed",
  1881 => x"4d2687c4",
  1882 => x"4b264c26",
  1883 => x"5e0e4f26",
  1884 => x"0e5d5c5b",
  1885 => x"f3c24a71",
  1886 => x"724cbfe9",
  1887 => x"87cb029a",
  1888 => x"c191c849",
  1889 => x"714bccf4",
  1890 => x"c187c483",
  1891 => x"c04bccf8",
  1892 => x"7449134d",
  1893 => x"e5f3c299",
  1894 => x"d4ffb9bf",
  1895 => x"c1787148",
  1896 => x"c8852cb7",
  1897 => x"e804adb7",
  1898 => x"e1f3c287",
  1899 => x"80c848bf",
  1900 => x"58e5f3c2",
  1901 => x"1e87effe",
  1902 => x"4b711e73",
  1903 => x"029a4a13",
  1904 => x"497287cb",
  1905 => x"1387e7fe",
  1906 => x"f5059a4a",
  1907 => x"87dafe87",
  1908 => x"e1f3c21e",
  1909 => x"f3c249bf",
  1910 => x"a1c148e1",
  1911 => x"b7c0c478",
  1912 => x"87db03a9",
  1913 => x"c248d4ff",
  1914 => x"78bfe5f3",
  1915 => x"bfe1f3c2",
  1916 => x"e1f3c249",
  1917 => x"78a1c148",
  1918 => x"a9b7c0c4",
  1919 => x"ff87e504",
  1920 => x"78c848d0",
  1921 => x"48edf3c2",
  1922 => x"4f2678c0",
  1923 => x"00000000",
  1924 => x"00000000",
  1925 => x"5f000000",
  1926 => x"0000005f",
  1927 => x"00030300",
  1928 => x"00000303",
  1929 => x"147f7f14",
  1930 => x"00147f7f",
  1931 => x"6b2e2400",
  1932 => x"00123a6b",
  1933 => x"18366a4c",
  1934 => x"0032566c",
  1935 => x"594f7e30",
  1936 => x"40683a77",
  1937 => x"07040000",
  1938 => x"00000003",
  1939 => x"3e1c0000",
  1940 => x"00004163",
  1941 => x"63410000",
  1942 => x"00001c3e",
  1943 => x"1c3e2a08",
  1944 => x"082a3e1c",
  1945 => x"3e080800",
  1946 => x"0008083e",
  1947 => x"e0800000",
  1948 => x"00000060",
  1949 => x"08080800",
  1950 => x"00080808",
  1951 => x"60000000",
  1952 => x"00000060",
  1953 => x"18306040",
  1954 => x"0103060c",
  1955 => x"597f3e00",
  1956 => x"003e7f4d",
  1957 => x"7f060400",
  1958 => x"0000007f",
  1959 => x"71634200",
  1960 => x"00464f59",
  1961 => x"49632200",
  1962 => x"00367f49",
  1963 => x"13161c18",
  1964 => x"00107f7f",
  1965 => x"45672700",
  1966 => x"00397d45",
  1967 => x"4b7e3c00",
  1968 => x"00307949",
  1969 => x"71010100",
  1970 => x"00070f79",
  1971 => x"497f3600",
  1972 => x"00367f49",
  1973 => x"494f0600",
  1974 => x"001e3f69",
  1975 => x"66000000",
  1976 => x"00000066",
  1977 => x"e6800000",
  1978 => x"00000066",
  1979 => x"14080800",
  1980 => x"00222214",
  1981 => x"14141400",
  1982 => x"00141414",
  1983 => x"14222200",
  1984 => x"00080814",
  1985 => x"51030200",
  1986 => x"00060f59",
  1987 => x"5d417f3e",
  1988 => x"001e1f55",
  1989 => x"097f7e00",
  1990 => x"007e7f09",
  1991 => x"497f7f00",
  1992 => x"00367f49",
  1993 => x"633e1c00",
  1994 => x"00414141",
  1995 => x"417f7f00",
  1996 => x"001c3e63",
  1997 => x"497f7f00",
  1998 => x"00414149",
  1999 => x"097f7f00",
  2000 => x"00010109",
  2001 => x"417f3e00",
  2002 => x"007a7b49",
  2003 => x"087f7f00",
  2004 => x"007f7f08",
  2005 => x"7f410000",
  2006 => x"0000417f",
  2007 => x"40602000",
  2008 => x"003f7f40",
  2009 => x"1c087f7f",
  2010 => x"00416336",
  2011 => x"407f7f00",
  2012 => x"00404040",
  2013 => x"0c067f7f",
  2014 => x"007f7f06",
  2015 => x"0c067f7f",
  2016 => x"007f7f18",
  2017 => x"417f3e00",
  2018 => x"003e7f41",
  2019 => x"097f7f00",
  2020 => x"00060f09",
  2021 => x"61417f3e",
  2022 => x"00407e7f",
  2023 => x"097f7f00",
  2024 => x"00667f19",
  2025 => x"4d6f2600",
  2026 => x"00327b59",
  2027 => x"7f010100",
  2028 => x"0001017f",
  2029 => x"407f3f00",
  2030 => x"003f7f40",
  2031 => x"703f0f00",
  2032 => x"000f3f70",
  2033 => x"18307f7f",
  2034 => x"007f7f30",
  2035 => x"1c366341",
  2036 => x"4163361c",
  2037 => x"7c060301",
  2038 => x"0103067c",
  2039 => x"4d597161",
  2040 => x"00414347",
  2041 => x"7f7f0000",
  2042 => x"00004141",
  2043 => x"0c060301",
  2044 => x"40603018",
  2045 => x"41410000",
  2046 => x"00007f7f",
  2047 => x"03060c08",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
