
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f0",x"f6",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"f0",x"f6",x"c2"),
    14 => (x"48",x"d0",x"e2",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"ee",x"e1"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"11",x"1e",x"4f"),
    50 => (x"78",x"08",x"d4",x"ff"),
    51 => (x"c1",x"48",x"66",x"c4"),
    52 => (x"58",x"a6",x"c8",x"88"),
    53 => (x"ed",x"05",x"98",x"70"),
    54 => (x"1e",x"4f",x"26",x"87"),
    55 => (x"c3",x"48",x"d4",x"ff"),
    56 => (x"51",x"68",x"78",x"ff"),
    57 => (x"c1",x"48",x"66",x"c4"),
    58 => (x"58",x"a6",x"c8",x"88"),
    59 => (x"eb",x"05",x"98",x"70"),
    60 => (x"1e",x"4f",x"26",x"87"),
    61 => (x"d4",x"ff",x"1e",x"73"),
    62 => (x"7b",x"ff",x"c3",x"4b"),
    63 => (x"ff",x"c3",x"4a",x"6b"),
    64 => (x"c8",x"49",x"6b",x"7b"),
    65 => (x"c3",x"b1",x"72",x"32"),
    66 => (x"4a",x"6b",x"7b",x"ff"),
    67 => (x"b2",x"71",x"31",x"c8"),
    68 => (x"6b",x"7b",x"ff",x"c3"),
    69 => (x"72",x"32",x"c8",x"49"),
    70 => (x"c4",x"48",x"71",x"b1"),
    71 => (x"26",x"4d",x"26",x"87"),
    72 => (x"26",x"4b",x"26",x"4c"),
    73 => (x"5b",x"5e",x"0e",x"4f"),
    74 => (x"71",x"0e",x"5d",x"5c"),
    75 => (x"4c",x"d4",x"ff",x"4a"),
    76 => (x"ff",x"c3",x"49",x"72"),
    77 => (x"c2",x"7c",x"71",x"99"),
    78 => (x"05",x"bf",x"d0",x"e2"),
    79 => (x"66",x"d0",x"87",x"c8"),
    80 => (x"d4",x"30",x"c9",x"48"),
    81 => (x"66",x"d0",x"58",x"a6"),
    82 => (x"c3",x"29",x"d8",x"49"),
    83 => (x"7c",x"71",x"99",x"ff"),
    84 => (x"d0",x"49",x"66",x"d0"),
    85 => (x"99",x"ff",x"c3",x"29"),
    86 => (x"66",x"d0",x"7c",x"71"),
    87 => (x"c3",x"29",x"c8",x"49"),
    88 => (x"7c",x"71",x"99",x"ff"),
    89 => (x"c3",x"49",x"66",x"d0"),
    90 => (x"7c",x"71",x"99",x"ff"),
    91 => (x"29",x"d0",x"49",x"72"),
    92 => (x"71",x"99",x"ff",x"c3"),
    93 => (x"c9",x"4b",x"6c",x"7c"),
    94 => (x"c3",x"4d",x"ff",x"f0"),
    95 => (x"d0",x"05",x"ab",x"ff"),
    96 => (x"7c",x"ff",x"c3",x"87"),
    97 => (x"8d",x"c1",x"4b",x"6c"),
    98 => (x"c3",x"87",x"c6",x"02"),
    99 => (x"f0",x"02",x"ab",x"ff"),
   100 => (x"fe",x"48",x"73",x"87"),
   101 => (x"c0",x"1e",x"87",x"c7"),
   102 => (x"48",x"d4",x"ff",x"49"),
   103 => (x"c1",x"78",x"ff",x"c3"),
   104 => (x"b7",x"c8",x"c3",x"81"),
   105 => (x"87",x"f1",x"04",x"a9"),
   106 => (x"73",x"1e",x"4f",x"26"),
   107 => (x"c4",x"87",x"e7",x"1e"),
   108 => (x"c0",x"4b",x"df",x"f8"),
   109 => (x"f0",x"ff",x"c0",x"1e"),
   110 => (x"fd",x"49",x"f7",x"c1"),
   111 => (x"86",x"c4",x"87",x"e7"),
   112 => (x"c0",x"05",x"a8",x"c1"),
   113 => (x"d4",x"ff",x"87",x"ea"),
   114 => (x"78",x"ff",x"c3",x"48"),
   115 => (x"c0",x"c0",x"c0",x"c1"),
   116 => (x"c0",x"1e",x"c0",x"c0"),
   117 => (x"e9",x"c1",x"f0",x"e1"),
   118 => (x"87",x"c9",x"fd",x"49"),
   119 => (x"98",x"70",x"86",x"c4"),
   120 => (x"ff",x"87",x"ca",x"05"),
   121 => (x"ff",x"c3",x"48",x"d4"),
   122 => (x"cb",x"48",x"c1",x"78"),
   123 => (x"87",x"e6",x"fe",x"87"),
   124 => (x"fe",x"05",x"8b",x"c1"),
   125 => (x"48",x"c0",x"87",x"fd"),
   126 => (x"1e",x"87",x"e6",x"fc"),
   127 => (x"d4",x"ff",x"1e",x"73"),
   128 => (x"78",x"ff",x"c3",x"48"),
   129 => (x"1e",x"c0",x"4b",x"d3"),
   130 => (x"c1",x"f0",x"ff",x"c0"),
   131 => (x"d4",x"fc",x"49",x"c1"),
   132 => (x"70",x"86",x"c4",x"87"),
   133 => (x"87",x"ca",x"05",x"98"),
   134 => (x"c3",x"48",x"d4",x"ff"),
   135 => (x"48",x"c1",x"78",x"ff"),
   136 => (x"f1",x"fd",x"87",x"cb"),
   137 => (x"05",x"8b",x"c1",x"87"),
   138 => (x"c0",x"87",x"db",x"ff"),
   139 => (x"87",x"f1",x"fb",x"48"),
   140 => (x"5c",x"5b",x"5e",x"0e"),
   141 => (x"4c",x"d4",x"ff",x"0e"),
   142 => (x"c6",x"87",x"db",x"fd"),
   143 => (x"e1",x"c0",x"1e",x"ea"),
   144 => (x"49",x"c8",x"c1",x"f0"),
   145 => (x"c4",x"87",x"de",x"fb"),
   146 => (x"02",x"a8",x"c1",x"86"),
   147 => (x"ea",x"fe",x"87",x"c8"),
   148 => (x"c1",x"48",x"c0",x"87"),
   149 => (x"da",x"fa",x"87",x"e2"),
   150 => (x"cf",x"49",x"70",x"87"),
   151 => (x"c6",x"99",x"ff",x"ff"),
   152 => (x"c8",x"02",x"a9",x"ea"),
   153 => (x"87",x"d3",x"fe",x"87"),
   154 => (x"cb",x"c1",x"48",x"c0"),
   155 => (x"7c",x"ff",x"c3",x"87"),
   156 => (x"fc",x"4b",x"f1",x"c0"),
   157 => (x"98",x"70",x"87",x"f4"),
   158 => (x"87",x"eb",x"c0",x"02"),
   159 => (x"ff",x"c0",x"1e",x"c0"),
   160 => (x"49",x"fa",x"c1",x"f0"),
   161 => (x"c4",x"87",x"de",x"fa"),
   162 => (x"05",x"98",x"70",x"86"),
   163 => (x"ff",x"c3",x"87",x"d9"),
   164 => (x"c3",x"49",x"6c",x"7c"),
   165 => (x"7c",x"7c",x"7c",x"ff"),
   166 => (x"99",x"c0",x"c1",x"7c"),
   167 => (x"c1",x"87",x"c4",x"02"),
   168 => (x"c0",x"87",x"d5",x"48"),
   169 => (x"c2",x"87",x"d1",x"48"),
   170 => (x"87",x"c4",x"05",x"ab"),
   171 => (x"87",x"c8",x"48",x"c0"),
   172 => (x"fe",x"05",x"8b",x"c1"),
   173 => (x"48",x"c0",x"87",x"fd"),
   174 => (x"1e",x"87",x"e4",x"f9"),
   175 => (x"e2",x"c2",x"1e",x"73"),
   176 => (x"78",x"c1",x"48",x"d0"),
   177 => (x"d0",x"ff",x"4b",x"c7"),
   178 => (x"fb",x"78",x"c2",x"48"),
   179 => (x"d0",x"ff",x"87",x"c8"),
   180 => (x"c0",x"78",x"c3",x"48"),
   181 => (x"d0",x"e5",x"c0",x"1e"),
   182 => (x"f9",x"49",x"c0",x"c1"),
   183 => (x"86",x"c4",x"87",x"c7"),
   184 => (x"c1",x"05",x"a8",x"c1"),
   185 => (x"ab",x"c2",x"4b",x"87"),
   186 => (x"c0",x"87",x"c5",x"05"),
   187 => (x"87",x"f9",x"c0",x"48"),
   188 => (x"ff",x"05",x"8b",x"c1"),
   189 => (x"f7",x"fc",x"87",x"d0"),
   190 => (x"d4",x"e2",x"c2",x"87"),
   191 => (x"05",x"98",x"70",x"58"),
   192 => (x"1e",x"c1",x"87",x"cd"),
   193 => (x"c1",x"f0",x"ff",x"c0"),
   194 => (x"d8",x"f8",x"49",x"d0"),
   195 => (x"ff",x"86",x"c4",x"87"),
   196 => (x"ff",x"c3",x"48",x"d4"),
   197 => (x"87",x"e0",x"c4",x"78"),
   198 => (x"58",x"d8",x"e2",x"c2"),
   199 => (x"c2",x"48",x"d0",x"ff"),
   200 => (x"48",x"d4",x"ff",x"78"),
   201 => (x"c1",x"78",x"ff",x"c3"),
   202 => (x"87",x"f5",x"f7",x"48"),
   203 => (x"5c",x"5b",x"5e",x"0e"),
   204 => (x"4a",x"71",x"0e",x"5d"),
   205 => (x"ff",x"4d",x"ff",x"c3"),
   206 => (x"7c",x"75",x"4c",x"d4"),
   207 => (x"c4",x"48",x"d0",x"ff"),
   208 => (x"7c",x"75",x"78",x"c3"),
   209 => (x"ff",x"c0",x"1e",x"72"),
   210 => (x"49",x"d8",x"c1",x"f0"),
   211 => (x"c4",x"87",x"d6",x"f7"),
   212 => (x"02",x"98",x"70",x"86"),
   213 => (x"48",x"c0",x"87",x"c5"),
   214 => (x"75",x"87",x"f0",x"c0"),
   215 => (x"7c",x"fe",x"c3",x"7c"),
   216 => (x"d4",x"1e",x"c0",x"c8"),
   217 => (x"dc",x"f5",x"49",x"66"),
   218 => (x"75",x"86",x"c4",x"87"),
   219 => (x"75",x"7c",x"75",x"7c"),
   220 => (x"e0",x"da",x"d8",x"7c"),
   221 => (x"6c",x"7c",x"75",x"4b"),
   222 => (x"c5",x"05",x"99",x"49"),
   223 => (x"05",x"8b",x"c1",x"87"),
   224 => (x"7c",x"75",x"87",x"f3"),
   225 => (x"c2",x"48",x"d0",x"ff"),
   226 => (x"f6",x"48",x"c1",x"78"),
   227 => (x"ff",x"1e",x"87",x"cf"),
   228 => (x"d0",x"ff",x"4a",x"d4"),
   229 => (x"78",x"d1",x"c4",x"48"),
   230 => (x"c1",x"7a",x"ff",x"c3"),
   231 => (x"87",x"f8",x"05",x"89"),
   232 => (x"73",x"1e",x"4f",x"26"),
   233 => (x"c5",x"4b",x"71",x"1e"),
   234 => (x"4a",x"df",x"cd",x"ee"),
   235 => (x"c3",x"48",x"d4",x"ff"),
   236 => (x"48",x"68",x"78",x"ff"),
   237 => (x"02",x"a8",x"fe",x"c3"),
   238 => (x"8a",x"c1",x"87",x"c5"),
   239 => (x"72",x"87",x"ed",x"05"),
   240 => (x"87",x"c5",x"05",x"9a"),
   241 => (x"ea",x"c0",x"48",x"c0"),
   242 => (x"02",x"9b",x"73",x"87"),
   243 => (x"66",x"c8",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c5"),
   246 => (x"66",x"c8",x"87",x"c6"),
   247 => (x"87",x"ee",x"fe",x"49"),
   248 => (x"c3",x"48",x"d4",x"ff"),
   249 => (x"73",x"78",x"78",x"ff"),
   250 => (x"87",x"c5",x"05",x"9b"),
   251 => (x"d0",x"48",x"d0",x"ff"),
   252 => (x"f4",x"48",x"c1",x"78"),
   253 => (x"73",x"1e",x"87",x"eb"),
   254 => (x"c0",x"4a",x"71",x"1e"),
   255 => (x"48",x"d4",x"ff",x"4b"),
   256 => (x"ff",x"78",x"ff",x"c3"),
   257 => (x"c3",x"c4",x"48",x"d0"),
   258 => (x"48",x"d4",x"ff",x"78"),
   259 => (x"72",x"78",x"ff",x"c3"),
   260 => (x"f0",x"ff",x"c0",x"1e"),
   261 => (x"f4",x"49",x"d1",x"c1"),
   262 => (x"86",x"c4",x"87",x"cb"),
   263 => (x"cd",x"05",x"98",x"70"),
   264 => (x"1e",x"c0",x"c8",x"87"),
   265 => (x"fd",x"49",x"66",x"cc"),
   266 => (x"86",x"c4",x"87",x"f8"),
   267 => (x"d0",x"ff",x"4b",x"70"),
   268 => (x"73",x"78",x"c2",x"48"),
   269 => (x"87",x"e9",x"f3",x"48"),
   270 => (x"5c",x"5b",x"5e",x"0e"),
   271 => (x"1e",x"c0",x"0e",x"5d"),
   272 => (x"c1",x"f0",x"ff",x"c0"),
   273 => (x"dc",x"f3",x"49",x"c9"),
   274 => (x"c2",x"1e",x"d2",x"87"),
   275 => (x"fd",x"49",x"d8",x"e2"),
   276 => (x"86",x"c8",x"87",x"d0"),
   277 => (x"84",x"c1",x"4c",x"c0"),
   278 => (x"04",x"ac",x"b7",x"d2"),
   279 => (x"e2",x"c2",x"87",x"f8"),
   280 => (x"49",x"bf",x"97",x"d8"),
   281 => (x"c1",x"99",x"c0",x"c3"),
   282 => (x"c0",x"05",x"a9",x"c0"),
   283 => (x"e2",x"c2",x"87",x"e7"),
   284 => (x"49",x"bf",x"97",x"df"),
   285 => (x"e2",x"c2",x"31",x"d0"),
   286 => (x"4a",x"bf",x"97",x"e0"),
   287 => (x"b1",x"72",x"32",x"c8"),
   288 => (x"97",x"e1",x"e2",x"c2"),
   289 => (x"71",x"b1",x"4a",x"bf"),
   290 => (x"ff",x"ff",x"cf",x"4c"),
   291 => (x"84",x"c1",x"9c",x"ff"),
   292 => (x"e7",x"c1",x"34",x"ca"),
   293 => (x"e1",x"e2",x"c2",x"87"),
   294 => (x"c1",x"49",x"bf",x"97"),
   295 => (x"c2",x"99",x"c6",x"31"),
   296 => (x"bf",x"97",x"e2",x"e2"),
   297 => (x"2a",x"b7",x"c7",x"4a"),
   298 => (x"e2",x"c2",x"b1",x"72"),
   299 => (x"4a",x"bf",x"97",x"dd"),
   300 => (x"c2",x"9d",x"cf",x"4d"),
   301 => (x"bf",x"97",x"de",x"e2"),
   302 => (x"ca",x"9a",x"c3",x"4a"),
   303 => (x"df",x"e2",x"c2",x"32"),
   304 => (x"c2",x"4b",x"bf",x"97"),
   305 => (x"c2",x"b2",x"73",x"33"),
   306 => (x"bf",x"97",x"e0",x"e2"),
   307 => (x"9b",x"c0",x"c3",x"4b"),
   308 => (x"73",x"2b",x"b7",x"c6"),
   309 => (x"c1",x"81",x"c2",x"b2"),
   310 => (x"70",x"30",x"71",x"48"),
   311 => (x"75",x"48",x"c1",x"49"),
   312 => (x"72",x"4d",x"70",x"30"),
   313 => (x"71",x"84",x"c1",x"4c"),
   314 => (x"b7",x"c0",x"c8",x"94"),
   315 => (x"87",x"cc",x"06",x"ad"),
   316 => (x"2d",x"b7",x"34",x"c1"),
   317 => (x"ad",x"b7",x"c0",x"c8"),
   318 => (x"87",x"f4",x"ff",x"01"),
   319 => (x"dc",x"f0",x"48",x"74"),
   320 => (x"5b",x"5e",x"0e",x"87"),
   321 => (x"f8",x"0e",x"5d",x"5c"),
   322 => (x"fe",x"ea",x"c2",x"86"),
   323 => (x"c2",x"78",x"c0",x"48"),
   324 => (x"c0",x"1e",x"f6",x"e2"),
   325 => (x"87",x"de",x"fb",x"49"),
   326 => (x"98",x"70",x"86",x"c4"),
   327 => (x"c0",x"87",x"c5",x"05"),
   328 => (x"87",x"ce",x"c9",x"48"),
   329 => (x"7e",x"c1",x"4d",x"c0"),
   330 => (x"bf",x"d0",x"f8",x"c0"),
   331 => (x"ec",x"e3",x"c2",x"49"),
   332 => (x"4b",x"c8",x"71",x"4a"),
   333 => (x"70",x"87",x"f3",x"ec"),
   334 => (x"87",x"c2",x"05",x"98"),
   335 => (x"f8",x"c0",x"7e",x"c0"),
   336 => (x"c2",x"49",x"bf",x"cc"),
   337 => (x"71",x"4a",x"c8",x"e4"),
   338 => (x"dd",x"ec",x"4b",x"c8"),
   339 => (x"05",x"98",x"70",x"87"),
   340 => (x"7e",x"c0",x"87",x"c2"),
   341 => (x"fd",x"c0",x"02",x"6e"),
   342 => (x"fc",x"e9",x"c2",x"87"),
   343 => (x"ea",x"c2",x"4d",x"bf"),
   344 => (x"7e",x"bf",x"9f",x"f4"),
   345 => (x"ea",x"d6",x"c5",x"48"),
   346 => (x"87",x"c7",x"05",x"a8"),
   347 => (x"bf",x"fc",x"e9",x"c2"),
   348 => (x"6e",x"87",x"ce",x"4d"),
   349 => (x"d5",x"e9",x"ca",x"48"),
   350 => (x"87",x"c5",x"02",x"a8"),
   351 => (x"f1",x"c7",x"48",x"c0"),
   352 => (x"f6",x"e2",x"c2",x"87"),
   353 => (x"f9",x"49",x"75",x"1e"),
   354 => (x"86",x"c4",x"87",x"ec"),
   355 => (x"c5",x"05",x"98",x"70"),
   356 => (x"c7",x"48",x"c0",x"87"),
   357 => (x"f8",x"c0",x"87",x"dc"),
   358 => (x"c2",x"49",x"bf",x"cc"),
   359 => (x"71",x"4a",x"c8",x"e4"),
   360 => (x"c5",x"eb",x"4b",x"c8"),
   361 => (x"05",x"98",x"70",x"87"),
   362 => (x"ea",x"c2",x"87",x"c8"),
   363 => (x"78",x"c1",x"48",x"fe"),
   364 => (x"f8",x"c0",x"87",x"da"),
   365 => (x"c2",x"49",x"bf",x"d0"),
   366 => (x"71",x"4a",x"ec",x"e3"),
   367 => (x"e9",x"ea",x"4b",x"c8"),
   368 => (x"02",x"98",x"70",x"87"),
   369 => (x"c0",x"87",x"c5",x"c0"),
   370 => (x"87",x"e6",x"c6",x"48"),
   371 => (x"97",x"f4",x"ea",x"c2"),
   372 => (x"d5",x"c1",x"49",x"bf"),
   373 => (x"cd",x"c0",x"05",x"a9"),
   374 => (x"f5",x"ea",x"c2",x"87"),
   375 => (x"c2",x"49",x"bf",x"97"),
   376 => (x"c0",x"02",x"a9",x"ea"),
   377 => (x"48",x"c0",x"87",x"c5"),
   378 => (x"c2",x"87",x"c7",x"c6"),
   379 => (x"bf",x"97",x"f6",x"e2"),
   380 => (x"e9",x"c3",x"48",x"7e"),
   381 => (x"ce",x"c0",x"02",x"a8"),
   382 => (x"c3",x"48",x"6e",x"87"),
   383 => (x"c0",x"02",x"a8",x"eb"),
   384 => (x"48",x"c0",x"87",x"c5"),
   385 => (x"c2",x"87",x"eb",x"c5"),
   386 => (x"bf",x"97",x"c1",x"e3"),
   387 => (x"c0",x"05",x"99",x"49"),
   388 => (x"e3",x"c2",x"87",x"cc"),
   389 => (x"49",x"bf",x"97",x"c2"),
   390 => (x"c0",x"02",x"a9",x"c2"),
   391 => (x"48",x"c0",x"87",x"c5"),
   392 => (x"c2",x"87",x"cf",x"c5"),
   393 => (x"bf",x"97",x"c3",x"e3"),
   394 => (x"fa",x"ea",x"c2",x"48"),
   395 => (x"48",x"4c",x"70",x"58"),
   396 => (x"ea",x"c2",x"88",x"c1"),
   397 => (x"e3",x"c2",x"58",x"fe"),
   398 => (x"49",x"bf",x"97",x"c4"),
   399 => (x"e3",x"c2",x"81",x"75"),
   400 => (x"4a",x"bf",x"97",x"c5"),
   401 => (x"a1",x"72",x"32",x"c8"),
   402 => (x"cb",x"ef",x"c2",x"7e"),
   403 => (x"c2",x"78",x"6e",x"48"),
   404 => (x"bf",x"97",x"c6",x"e3"),
   405 => (x"58",x"a6",x"c8",x"48"),
   406 => (x"bf",x"fe",x"ea",x"c2"),
   407 => (x"87",x"d4",x"c2",x"02"),
   408 => (x"bf",x"cc",x"f8",x"c0"),
   409 => (x"c8",x"e4",x"c2",x"49"),
   410 => (x"4b",x"c8",x"71",x"4a"),
   411 => (x"70",x"87",x"fb",x"e7"),
   412 => (x"c5",x"c0",x"02",x"98"),
   413 => (x"c3",x"48",x"c0",x"87"),
   414 => (x"ea",x"c2",x"87",x"f8"),
   415 => (x"c2",x"4c",x"bf",x"f6"),
   416 => (x"c2",x"5c",x"df",x"ef"),
   417 => (x"bf",x"97",x"db",x"e3"),
   418 => (x"c2",x"31",x"c8",x"49"),
   419 => (x"bf",x"97",x"da",x"e3"),
   420 => (x"c2",x"49",x"a1",x"4a"),
   421 => (x"bf",x"97",x"dc",x"e3"),
   422 => (x"72",x"32",x"d0",x"4a"),
   423 => (x"e3",x"c2",x"49",x"a1"),
   424 => (x"4a",x"bf",x"97",x"dd"),
   425 => (x"a1",x"72",x"32",x"d8"),
   426 => (x"91",x"66",x"c4",x"49"),
   427 => (x"bf",x"cb",x"ef",x"c2"),
   428 => (x"d3",x"ef",x"c2",x"81"),
   429 => (x"e3",x"e3",x"c2",x"59"),
   430 => (x"c8",x"4a",x"bf",x"97"),
   431 => (x"e2",x"e3",x"c2",x"32"),
   432 => (x"a2",x"4b",x"bf",x"97"),
   433 => (x"e4",x"e3",x"c2",x"4a"),
   434 => (x"d0",x"4b",x"bf",x"97"),
   435 => (x"4a",x"a2",x"73",x"33"),
   436 => (x"97",x"e5",x"e3",x"c2"),
   437 => (x"9b",x"cf",x"4b",x"bf"),
   438 => (x"a2",x"73",x"33",x"d8"),
   439 => (x"d7",x"ef",x"c2",x"4a"),
   440 => (x"d3",x"ef",x"c2",x"5a"),
   441 => (x"8a",x"c2",x"4a",x"bf"),
   442 => (x"ef",x"c2",x"92",x"74"),
   443 => (x"a1",x"72",x"48",x"d7"),
   444 => (x"87",x"ca",x"c1",x"78"),
   445 => (x"97",x"c8",x"e3",x"c2"),
   446 => (x"31",x"c8",x"49",x"bf"),
   447 => (x"97",x"c7",x"e3",x"c2"),
   448 => (x"49",x"a1",x"4a",x"bf"),
   449 => (x"59",x"c6",x"eb",x"c2"),
   450 => (x"bf",x"c2",x"eb",x"c2"),
   451 => (x"c7",x"31",x"c5",x"49"),
   452 => (x"29",x"c9",x"81",x"ff"),
   453 => (x"59",x"df",x"ef",x"c2"),
   454 => (x"97",x"cd",x"e3",x"c2"),
   455 => (x"32",x"c8",x"4a",x"bf"),
   456 => (x"97",x"cc",x"e3",x"c2"),
   457 => (x"4a",x"a2",x"4b",x"bf"),
   458 => (x"6e",x"92",x"66",x"c4"),
   459 => (x"db",x"ef",x"c2",x"82"),
   460 => (x"d3",x"ef",x"c2",x"5a"),
   461 => (x"c2",x"78",x"c0",x"48"),
   462 => (x"72",x"48",x"cf",x"ef"),
   463 => (x"ef",x"c2",x"78",x"a1"),
   464 => (x"ef",x"c2",x"48",x"df"),
   465 => (x"c2",x"78",x"bf",x"d3"),
   466 => (x"c2",x"48",x"e3",x"ef"),
   467 => (x"78",x"bf",x"d7",x"ef"),
   468 => (x"bf",x"fe",x"ea",x"c2"),
   469 => (x"87",x"c9",x"c0",x"02"),
   470 => (x"30",x"c4",x"48",x"74"),
   471 => (x"c9",x"c0",x"7e",x"70"),
   472 => (x"db",x"ef",x"c2",x"87"),
   473 => (x"30",x"c4",x"48",x"bf"),
   474 => (x"eb",x"c2",x"7e",x"70"),
   475 => (x"78",x"6e",x"48",x"c2"),
   476 => (x"8e",x"f8",x"48",x"c1"),
   477 => (x"4c",x"26",x"4d",x"26"),
   478 => (x"4f",x"26",x"4b",x"26"),
   479 => (x"5c",x"5b",x"5e",x"0e"),
   480 => (x"4a",x"71",x"0e",x"5d"),
   481 => (x"bf",x"fe",x"ea",x"c2"),
   482 => (x"72",x"87",x"cb",x"02"),
   483 => (x"72",x"2b",x"c7",x"4b"),
   484 => (x"9c",x"ff",x"c1",x"4c"),
   485 => (x"4b",x"72",x"87",x"c9"),
   486 => (x"4c",x"72",x"2b",x"c8"),
   487 => (x"c2",x"9c",x"ff",x"c3"),
   488 => (x"83",x"bf",x"cb",x"ef"),
   489 => (x"bf",x"c8",x"f8",x"c0"),
   490 => (x"87",x"d9",x"02",x"ab"),
   491 => (x"5b",x"cc",x"f8",x"c0"),
   492 => (x"1e",x"f6",x"e2",x"c2"),
   493 => (x"fd",x"f0",x"49",x"73"),
   494 => (x"70",x"86",x"c4",x"87"),
   495 => (x"87",x"c5",x"05",x"98"),
   496 => (x"e6",x"c0",x"48",x"c0"),
   497 => (x"fe",x"ea",x"c2",x"87"),
   498 => (x"87",x"d2",x"02",x"bf"),
   499 => (x"91",x"c4",x"49",x"74"),
   500 => (x"81",x"f6",x"e2",x"c2"),
   501 => (x"ff",x"cf",x"4d",x"69"),
   502 => (x"9d",x"ff",x"ff",x"ff"),
   503 => (x"49",x"74",x"87",x"cb"),
   504 => (x"e2",x"c2",x"91",x"c2"),
   505 => (x"69",x"9f",x"81",x"f6"),
   506 => (x"fe",x"48",x"75",x"4d"),
   507 => (x"5e",x"0e",x"87",x"c6"),
   508 => (x"0e",x"5d",x"5c",x"5b"),
   509 => (x"c0",x"4d",x"71",x"1e"),
   510 => (x"d0",x"49",x"c1",x"1e"),
   511 => (x"86",x"c4",x"87",x"f2"),
   512 => (x"02",x"9c",x"4c",x"70"),
   513 => (x"c2",x"87",x"c0",x"c1"),
   514 => (x"75",x"4a",x"c6",x"eb"),
   515 => (x"87",x"ff",x"e0",x"49"),
   516 => (x"c0",x"02",x"98",x"70"),
   517 => (x"4a",x"74",x"87",x"f1"),
   518 => (x"4b",x"cb",x"49",x"75"),
   519 => (x"70",x"87",x"e5",x"e1"),
   520 => (x"e2",x"c0",x"02",x"98"),
   521 => (x"74",x"1e",x"c0",x"87"),
   522 => (x"87",x"c7",x"02",x"9c"),
   523 => (x"c0",x"48",x"a6",x"c4"),
   524 => (x"c4",x"87",x"c5",x"78"),
   525 => (x"78",x"c1",x"48",x"a6"),
   526 => (x"cf",x"49",x"66",x"c4"),
   527 => (x"86",x"c4",x"87",x"f2"),
   528 => (x"05",x"9c",x"4c",x"70"),
   529 => (x"74",x"87",x"c0",x"ff"),
   530 => (x"e7",x"fc",x"26",x"48"),
   531 => (x"5b",x"5e",x"0e",x"87"),
   532 => (x"f8",x"0e",x"5d",x"5c"),
   533 => (x"9b",x"4b",x"71",x"86"),
   534 => (x"c0",x"87",x"c5",x"05"),
   535 => (x"87",x"d4",x"c2",x"48"),
   536 => (x"c0",x"4d",x"a3",x"c8"),
   537 => (x"02",x"66",x"d8",x"7d"),
   538 => (x"66",x"d8",x"87",x"c7"),
   539 => (x"c5",x"05",x"bf",x"97"),
   540 => (x"c1",x"48",x"c0",x"87"),
   541 => (x"66",x"d8",x"87",x"fe"),
   542 => (x"87",x"f2",x"fd",x"49"),
   543 => (x"02",x"6e",x"7e",x"70"),
   544 => (x"6e",x"87",x"ef",x"c1"),
   545 => (x"69",x"81",x"dc",x"49"),
   546 => (x"da",x"49",x"6e",x"7d"),
   547 => (x"4c",x"a3",x"c4",x"81"),
   548 => (x"c2",x"7c",x"69",x"9f"),
   549 => (x"02",x"bf",x"fe",x"ea"),
   550 => (x"49",x"6e",x"87",x"d0"),
   551 => (x"69",x"9f",x"81",x"d4"),
   552 => (x"ff",x"c0",x"4a",x"49"),
   553 => (x"32",x"d0",x"9a",x"ff"),
   554 => (x"4a",x"c0",x"87",x"c2"),
   555 => (x"6c",x"48",x"49",x"72"),
   556 => (x"c0",x"7c",x"70",x"80"),
   557 => (x"49",x"a3",x"cc",x"7b"),
   558 => (x"a3",x"d0",x"79",x"6c"),
   559 => (x"c4",x"79",x"c0",x"49"),
   560 => (x"78",x"c0",x"48",x"a6"),
   561 => (x"c4",x"4a",x"a3",x"d4"),
   562 => (x"91",x"c8",x"49",x"66"),
   563 => (x"c0",x"49",x"a1",x"72"),
   564 => (x"c4",x"79",x"6c",x"41"),
   565 => (x"80",x"c1",x"48",x"66"),
   566 => (x"c4",x"58",x"a6",x"c8"),
   567 => (x"ff",x"04",x"a8",x"b7"),
   568 => (x"4a",x"6d",x"87",x"e2"),
   569 => (x"2a",x"c5",x"2a",x"c9"),
   570 => (x"49",x"a3",x"f4",x"c0"),
   571 => (x"48",x"6e",x"79",x"72"),
   572 => (x"48",x"c0",x"87",x"c2"),
   573 => (x"fb",x"f9",x"8e",x"f8"),
   574 => (x"5b",x"5e",x"0e",x"87"),
   575 => (x"71",x"0e",x"5d",x"5c"),
   576 => (x"c8",x"f8",x"c0",x"4c"),
   577 => (x"74",x"78",x"ff",x"48"),
   578 => (x"ca",x"c1",x"02",x"9c"),
   579 => (x"49",x"a4",x"c8",x"87"),
   580 => (x"c2",x"c1",x"02",x"69"),
   581 => (x"4a",x"66",x"d0",x"87"),
   582 => (x"d4",x"82",x"49",x"6c"),
   583 => (x"66",x"d0",x"5a",x"a6"),
   584 => (x"ea",x"c2",x"b9",x"4d"),
   585 => (x"ff",x"4a",x"bf",x"fa"),
   586 => (x"71",x"99",x"72",x"ba"),
   587 => (x"e4",x"c0",x"02",x"99"),
   588 => (x"4b",x"a4",x"c4",x"87"),
   589 => (x"c3",x"f9",x"49",x"6b"),
   590 => (x"c2",x"7b",x"70",x"87"),
   591 => (x"49",x"bf",x"f6",x"ea"),
   592 => (x"7c",x"71",x"81",x"6c"),
   593 => (x"ea",x"c2",x"b9",x"75"),
   594 => (x"ff",x"4a",x"bf",x"fa"),
   595 => (x"71",x"99",x"72",x"ba"),
   596 => (x"dc",x"ff",x"05",x"99"),
   597 => (x"f8",x"7c",x"75",x"87"),
   598 => (x"73",x"1e",x"87",x"da"),
   599 => (x"9b",x"4b",x"71",x"1e"),
   600 => (x"c8",x"87",x"c7",x"02"),
   601 => (x"05",x"69",x"49",x"a3"),
   602 => (x"48",x"c0",x"87",x"c5"),
   603 => (x"c2",x"87",x"eb",x"c0"),
   604 => (x"4a",x"bf",x"cf",x"ef"),
   605 => (x"69",x"49",x"a3",x"c4"),
   606 => (x"c2",x"89",x"c2",x"49"),
   607 => (x"91",x"bf",x"f6",x"ea"),
   608 => (x"c2",x"4a",x"a2",x"71"),
   609 => (x"49",x"bf",x"fa",x"ea"),
   610 => (x"a2",x"71",x"99",x"6b"),
   611 => (x"1e",x"66",x"c8",x"4a"),
   612 => (x"e1",x"e9",x"49",x"72"),
   613 => (x"70",x"86",x"c4",x"87"),
   614 => (x"db",x"f7",x"48",x"49"),
   615 => (x"1e",x"73",x"1e",x"87"),
   616 => (x"02",x"9b",x"4b",x"71"),
   617 => (x"a3",x"c8",x"87",x"c7"),
   618 => (x"c5",x"05",x"69",x"49"),
   619 => (x"c0",x"48",x"c0",x"87"),
   620 => (x"ef",x"c2",x"87",x"eb"),
   621 => (x"c4",x"4a",x"bf",x"cf"),
   622 => (x"49",x"69",x"49",x"a3"),
   623 => (x"ea",x"c2",x"89",x"c2"),
   624 => (x"71",x"91",x"bf",x"f6"),
   625 => (x"ea",x"c2",x"4a",x"a2"),
   626 => (x"6b",x"49",x"bf",x"fa"),
   627 => (x"4a",x"a2",x"71",x"99"),
   628 => (x"72",x"1e",x"66",x"c8"),
   629 => (x"87",x"d4",x"e5",x"49"),
   630 => (x"49",x"70",x"86",x"c4"),
   631 => (x"87",x"d8",x"f6",x"48"),
   632 => (x"5c",x"5b",x"5e",x"0e"),
   633 => (x"86",x"f8",x"0e",x"5d"),
   634 => (x"a6",x"c4",x"4b",x"71"),
   635 => (x"c8",x"78",x"ff",x"48"),
   636 => (x"4d",x"69",x"49",x"a3"),
   637 => (x"a3",x"d4",x"4c",x"c0"),
   638 => (x"c8",x"49",x"74",x"4a"),
   639 => (x"49",x"a1",x"72",x"91"),
   640 => (x"66",x"d8",x"49",x"69"),
   641 => (x"70",x"88",x"71",x"48"),
   642 => (x"a9",x"66",x"d8",x"7e"),
   643 => (x"6e",x"87",x"ca",x"01"),
   644 => (x"87",x"c5",x"06",x"ad"),
   645 => (x"6e",x"5c",x"a6",x"c8"),
   646 => (x"c4",x"84",x"c1",x"4d"),
   647 => (x"ff",x"04",x"ac",x"b7"),
   648 => (x"48",x"66",x"87",x"d4"),
   649 => (x"cb",x"f5",x"8e",x"f8"),
   650 => (x"5b",x"5e",x"0e",x"87"),
   651 => (x"ec",x"0e",x"5d",x"5c"),
   652 => (x"59",x"a6",x"c8",x"86"),
   653 => (x"c1",x"48",x"a6",x"c8"),
   654 => (x"ff",x"ff",x"ff",x"ff"),
   655 => (x"80",x"c4",x"78",x"ff"),
   656 => (x"4d",x"c0",x"78",x"ff"),
   657 => (x"66",x"c4",x"4c",x"c0"),
   658 => (x"74",x"83",x"d4",x"4b"),
   659 => (x"73",x"91",x"c8",x"49"),
   660 => (x"4a",x"75",x"49",x"a1"),
   661 => (x"a2",x"73",x"92",x"c8"),
   662 => (x"6e",x"49",x"69",x"7e"),
   663 => (x"a6",x"d4",x"89",x"bf"),
   664 => (x"05",x"ad",x"74",x"59"),
   665 => (x"a6",x"d0",x"87",x"c6"),
   666 => (x"78",x"bf",x"6e",x"48"),
   667 => (x"c0",x"48",x"66",x"d0"),
   668 => (x"cf",x"04",x"a8",x"b7"),
   669 => (x"49",x"66",x"d0",x"87"),
   670 => (x"03",x"a9",x"66",x"c8"),
   671 => (x"a6",x"d0",x"87",x"c6"),
   672 => (x"59",x"a6",x"cc",x"5c"),
   673 => (x"b7",x"c4",x"84",x"c1"),
   674 => (x"f9",x"fe",x"04",x"ac"),
   675 => (x"c4",x"85",x"c1",x"87"),
   676 => (x"fe",x"04",x"ad",x"b7"),
   677 => (x"66",x"cc",x"87",x"ee"),
   678 => (x"f3",x"8e",x"ec",x"48"),
   679 => (x"5e",x"0e",x"87",x"d6"),
   680 => (x"0e",x"5d",x"5c",x"5b"),
   681 => (x"4b",x"71",x"86",x"f0"),
   682 => (x"4c",x"66",x"e0",x"c0"),
   683 => (x"9b",x"73",x"2c",x"c9"),
   684 => (x"87",x"e1",x"c3",x"02"),
   685 => (x"69",x"49",x"a3",x"c8"),
   686 => (x"87",x"d9",x"c3",x"02"),
   687 => (x"c0",x"49",x"a3",x"d0"),
   688 => (x"6b",x"79",x"66",x"e0"),
   689 => (x"c3",x"02",x"ac",x"7e"),
   690 => (x"ea",x"c2",x"87",x"cb"),
   691 => (x"ff",x"49",x"bf",x"fa"),
   692 => (x"74",x"4a",x"71",x"b9"),
   693 => (x"6e",x"48",x"71",x"9a"),
   694 => (x"58",x"a6",x"cc",x"98"),
   695 => (x"c4",x"4d",x"a3",x"c4"),
   696 => (x"78",x"6d",x"48",x"a6"),
   697 => (x"05",x"aa",x"66",x"c8"),
   698 => (x"7b",x"74",x"87",x"c5"),
   699 => (x"72",x"87",x"d1",x"c2"),
   700 => (x"fb",x"49",x"73",x"1e"),
   701 => (x"86",x"c4",x"87",x"ea"),
   702 => (x"c0",x"48",x"7e",x"70"),
   703 => (x"d0",x"04",x"a8",x"b7"),
   704 => (x"4a",x"a3",x"d4",x"87"),
   705 => (x"91",x"c8",x"49",x"6e"),
   706 => (x"21",x"49",x"a1",x"72"),
   707 => (x"c7",x"7d",x"69",x"7b"),
   708 => (x"cc",x"7b",x"c0",x"87"),
   709 => (x"7d",x"69",x"49",x"a3"),
   710 => (x"73",x"1e",x"66",x"c8"),
   711 => (x"87",x"c0",x"fb",x"49"),
   712 => (x"7e",x"70",x"86",x"c4"),
   713 => (x"49",x"a3",x"f4",x"c0"),
   714 => (x"69",x"48",x"a6",x"cc"),
   715 => (x"48",x"66",x"c8",x"78"),
   716 => (x"06",x"a8",x"66",x"cc"),
   717 => (x"48",x"6e",x"87",x"c9"),
   718 => (x"04",x"a8",x"b7",x"c0"),
   719 => (x"6e",x"87",x"e0",x"c0"),
   720 => (x"a8",x"b7",x"c0",x"48"),
   721 => (x"87",x"ec",x"c0",x"04"),
   722 => (x"6e",x"4a",x"a3",x"d4"),
   723 => (x"72",x"91",x"c8",x"49"),
   724 => (x"66",x"c8",x"49",x"a1"),
   725 => (x"70",x"88",x"69",x"48"),
   726 => (x"a9",x"66",x"cc",x"49"),
   727 => (x"73",x"87",x"d5",x"06"),
   728 => (x"87",x"c5",x"fb",x"49"),
   729 => (x"a3",x"d4",x"49",x"70"),
   730 => (x"72",x"91",x"c8",x"4a"),
   731 => (x"66",x"c8",x"49",x"a1"),
   732 => (x"79",x"66",x"c4",x"41"),
   733 => (x"49",x"74",x"8c",x"6b"),
   734 => (x"f5",x"49",x"73",x"1e"),
   735 => (x"86",x"c4",x"87",x"fb"),
   736 => (x"49",x"66",x"e0",x"c0"),
   737 => (x"02",x"99",x"ff",x"c7"),
   738 => (x"e2",x"c2",x"87",x"cb"),
   739 => (x"49",x"73",x"1e",x"f6"),
   740 => (x"c4",x"87",x"c7",x"f7"),
   741 => (x"ef",x"8e",x"f0",x"86"),
   742 => (x"73",x"1e",x"87",x"da"),
   743 => (x"9b",x"4b",x"71",x"1e"),
   744 => (x"87",x"e4",x"c0",x"02"),
   745 => (x"5b",x"e3",x"ef",x"c2"),
   746 => (x"8a",x"c2",x"4a",x"73"),
   747 => (x"bf",x"f6",x"ea",x"c2"),
   748 => (x"ef",x"c2",x"92",x"49"),
   749 => (x"72",x"48",x"bf",x"cf"),
   750 => (x"e7",x"ef",x"c2",x"80"),
   751 => (x"c4",x"48",x"71",x"58"),
   752 => (x"c6",x"eb",x"c2",x"30"),
   753 => (x"87",x"ed",x"c0",x"58"),
   754 => (x"48",x"df",x"ef",x"c2"),
   755 => (x"bf",x"d3",x"ef",x"c2"),
   756 => (x"e3",x"ef",x"c2",x"78"),
   757 => (x"d7",x"ef",x"c2",x"48"),
   758 => (x"ea",x"c2",x"78",x"bf"),
   759 => (x"c9",x"02",x"bf",x"fe"),
   760 => (x"f6",x"ea",x"c2",x"87"),
   761 => (x"31",x"c4",x"49",x"bf"),
   762 => (x"ef",x"c2",x"87",x"c7"),
   763 => (x"c4",x"49",x"bf",x"db"),
   764 => (x"c6",x"eb",x"c2",x"31"),
   765 => (x"87",x"c0",x"ee",x"59"),
   766 => (x"5c",x"5b",x"5e",x"0e"),
   767 => (x"c0",x"4a",x"71",x"0e"),
   768 => (x"02",x"9a",x"72",x"4b"),
   769 => (x"da",x"87",x"e1",x"c0"),
   770 => (x"69",x"9f",x"49",x"a2"),
   771 => (x"fe",x"ea",x"c2",x"4b"),
   772 => (x"87",x"cf",x"02",x"bf"),
   773 => (x"9f",x"49",x"a2",x"d4"),
   774 => (x"c0",x"4c",x"49",x"69"),
   775 => (x"d0",x"9c",x"ff",x"ff"),
   776 => (x"c0",x"87",x"c2",x"34"),
   777 => (x"b3",x"49",x"74",x"4c"),
   778 => (x"ed",x"fd",x"49",x"73"),
   779 => (x"87",x"c6",x"ed",x"87"),
   780 => (x"5c",x"5b",x"5e",x"0e"),
   781 => (x"86",x"f4",x"0e",x"5d"),
   782 => (x"7e",x"c0",x"4a",x"71"),
   783 => (x"d8",x"02",x"9a",x"72"),
   784 => (x"f2",x"e2",x"c2",x"87"),
   785 => (x"c2",x"78",x"c0",x"48"),
   786 => (x"c2",x"48",x"ea",x"e2"),
   787 => (x"78",x"bf",x"e3",x"ef"),
   788 => (x"48",x"ee",x"e2",x"c2"),
   789 => (x"bf",x"df",x"ef",x"c2"),
   790 => (x"d3",x"eb",x"c2",x"78"),
   791 => (x"c2",x"50",x"c0",x"48"),
   792 => (x"49",x"bf",x"c2",x"eb"),
   793 => (x"bf",x"f2",x"e2",x"c2"),
   794 => (x"03",x"aa",x"71",x"4a"),
   795 => (x"72",x"87",x"c0",x"c4"),
   796 => (x"05",x"99",x"cf",x"49"),
   797 => (x"c2",x"87",x"e1",x"c0"),
   798 => (x"c2",x"1e",x"f6",x"e2"),
   799 => (x"49",x"bf",x"ea",x"e2"),
   800 => (x"48",x"ea",x"e2",x"c2"),
   801 => (x"71",x"78",x"a1",x"c1"),
   802 => (x"87",x"ea",x"dd",x"ff"),
   803 => (x"f8",x"c0",x"86",x"c4"),
   804 => (x"e2",x"c2",x"48",x"c4"),
   805 => (x"87",x"cc",x"78",x"f6"),
   806 => (x"bf",x"c4",x"f8",x"c0"),
   807 => (x"80",x"e0",x"c0",x"48"),
   808 => (x"58",x"c8",x"f8",x"c0"),
   809 => (x"bf",x"f2",x"e2",x"c2"),
   810 => (x"c2",x"80",x"c1",x"48"),
   811 => (x"27",x"58",x"f6",x"e2"),
   812 => (x"00",x"00",x"0e",x"04"),
   813 => (x"4d",x"bf",x"97",x"bf"),
   814 => (x"e2",x"c2",x"02",x"9d"),
   815 => (x"ad",x"e5",x"c3",x"87"),
   816 => (x"87",x"db",x"c2",x"02"),
   817 => (x"bf",x"c4",x"f8",x"c0"),
   818 => (x"49",x"a3",x"cb",x"4b"),
   819 => (x"ac",x"cf",x"4c",x"11"),
   820 => (x"87",x"d2",x"c1",x"05"),
   821 => (x"99",x"df",x"49",x"75"),
   822 => (x"91",x"cd",x"89",x"c1"),
   823 => (x"81",x"c6",x"eb",x"c2"),
   824 => (x"12",x"4a",x"a3",x"c1"),
   825 => (x"4a",x"a3",x"c3",x"51"),
   826 => (x"a3",x"c5",x"51",x"12"),
   827 => (x"c7",x"51",x"12",x"4a"),
   828 => (x"51",x"12",x"4a",x"a3"),
   829 => (x"12",x"4a",x"a3",x"c9"),
   830 => (x"4a",x"a3",x"ce",x"51"),
   831 => (x"a3",x"d0",x"51",x"12"),
   832 => (x"d2",x"51",x"12",x"4a"),
   833 => (x"51",x"12",x"4a",x"a3"),
   834 => (x"12",x"4a",x"a3",x"d4"),
   835 => (x"4a",x"a3",x"d6",x"51"),
   836 => (x"a3",x"d8",x"51",x"12"),
   837 => (x"dc",x"51",x"12",x"4a"),
   838 => (x"51",x"12",x"4a",x"a3"),
   839 => (x"12",x"4a",x"a3",x"de"),
   840 => (x"c0",x"7e",x"c1",x"51"),
   841 => (x"49",x"74",x"87",x"f9"),
   842 => (x"c0",x"05",x"99",x"c8"),
   843 => (x"49",x"74",x"87",x"ea"),
   844 => (x"d0",x"05",x"99",x"d0"),
   845 => (x"02",x"66",x"dc",x"87"),
   846 => (x"73",x"87",x"ca",x"c0"),
   847 => (x"0f",x"66",x"dc",x"49"),
   848 => (x"d3",x"02",x"98",x"70"),
   849 => (x"c0",x"05",x"6e",x"87"),
   850 => (x"eb",x"c2",x"87",x"c6"),
   851 => (x"50",x"c0",x"48",x"c6"),
   852 => (x"bf",x"c4",x"f8",x"c0"),
   853 => (x"87",x"e7",x"c2",x"48"),
   854 => (x"48",x"d3",x"eb",x"c2"),
   855 => (x"c2",x"7e",x"50",x"c0"),
   856 => (x"49",x"bf",x"c2",x"eb"),
   857 => (x"bf",x"f2",x"e2",x"c2"),
   858 => (x"04",x"aa",x"71",x"4a"),
   859 => (x"c2",x"87",x"c0",x"fc"),
   860 => (x"05",x"bf",x"e3",x"ef"),
   861 => (x"c2",x"87",x"c8",x"c0"),
   862 => (x"02",x"bf",x"fe",x"ea"),
   863 => (x"c0",x"87",x"fe",x"c1"),
   864 => (x"ff",x"48",x"c8",x"f8"),
   865 => (x"ee",x"e2",x"c2",x"78"),
   866 => (x"ef",x"e7",x"49",x"bf"),
   867 => (x"c2",x"49",x"70",x"87"),
   868 => (x"c4",x"59",x"f2",x"e2"),
   869 => (x"e2",x"c2",x"48",x"a6"),
   870 => (x"c2",x"78",x"bf",x"ee"),
   871 => (x"02",x"bf",x"fe",x"ea"),
   872 => (x"c4",x"87",x"d8",x"c0"),
   873 => (x"ff",x"cf",x"49",x"66"),
   874 => (x"99",x"f8",x"ff",x"ff"),
   875 => (x"c5",x"c0",x"02",x"a9"),
   876 => (x"c0",x"4d",x"c0",x"87"),
   877 => (x"4d",x"c1",x"87",x"e1"),
   878 => (x"c4",x"87",x"dc",x"c0"),
   879 => (x"ff",x"cf",x"49",x"66"),
   880 => (x"02",x"a9",x"99",x"f8"),
   881 => (x"c8",x"87",x"c8",x"c0"),
   882 => (x"78",x"c0",x"48",x"a6"),
   883 => (x"c8",x"87",x"c5",x"c0"),
   884 => (x"78",x"c1",x"48",x"a6"),
   885 => (x"75",x"4d",x"66",x"c8"),
   886 => (x"e0",x"c0",x"05",x"9d"),
   887 => (x"49",x"66",x"c4",x"87"),
   888 => (x"ea",x"c2",x"89",x"c2"),
   889 => (x"91",x"4a",x"bf",x"f6"),
   890 => (x"bf",x"cf",x"ef",x"c2"),
   891 => (x"ea",x"e2",x"c2",x"4a"),
   892 => (x"78",x"a1",x"72",x"48"),
   893 => (x"48",x"f2",x"e2",x"c2"),
   894 => (x"e2",x"f9",x"78",x"c0"),
   895 => (x"f4",x"48",x"c0",x"87"),
   896 => (x"87",x"f0",x"e5",x"8e"),
   897 => (x"00",x"00",x"00",x"00"),
   898 => (x"ff",x"ff",x"ff",x"ff"),
   899 => (x"00",x"00",x"0e",x"14"),
   900 => (x"00",x"00",x"0e",x"1d"),
   901 => (x"33",x"54",x"41",x"46"),
   902 => (x"20",x"20",x"20",x"32"),
   903 => (x"54",x"41",x"46",x"00"),
   904 => (x"20",x"20",x"36",x"31"),
   905 => (x"ff",x"1e",x"00",x"20"),
   906 => (x"ff",x"c3",x"48",x"d4"),
   907 => (x"26",x"48",x"68",x"78"),
   908 => (x"d4",x"ff",x"1e",x"4f"),
   909 => (x"78",x"ff",x"c3",x"48"),
   910 => (x"c8",x"48",x"d0",x"ff"),
   911 => (x"d4",x"ff",x"78",x"e1"),
   912 => (x"c2",x"78",x"d4",x"48"),
   913 => (x"ff",x"48",x"e7",x"ef"),
   914 => (x"26",x"50",x"bf",x"d4"),
   915 => (x"d0",x"ff",x"1e",x"4f"),
   916 => (x"78",x"e0",x"c0",x"48"),
   917 => (x"ff",x"1e",x"4f",x"26"),
   918 => (x"49",x"70",x"87",x"cc"),
   919 => (x"87",x"c6",x"02",x"99"),
   920 => (x"05",x"a9",x"fb",x"c0"),
   921 => (x"48",x"71",x"87",x"f1"),
   922 => (x"5e",x"0e",x"4f",x"26"),
   923 => (x"71",x"0e",x"5c",x"5b"),
   924 => (x"fe",x"4c",x"c0",x"4b"),
   925 => (x"49",x"70",x"87",x"f0"),
   926 => (x"f9",x"c0",x"02",x"99"),
   927 => (x"a9",x"ec",x"c0",x"87"),
   928 => (x"87",x"f2",x"c0",x"02"),
   929 => (x"02",x"a9",x"fb",x"c0"),
   930 => (x"cc",x"87",x"eb",x"c0"),
   931 => (x"03",x"ac",x"b7",x"66"),
   932 => (x"66",x"d0",x"87",x"c7"),
   933 => (x"71",x"87",x"c2",x"02"),
   934 => (x"02",x"99",x"71",x"53"),
   935 => (x"84",x"c1",x"87",x"c2"),
   936 => (x"70",x"87",x"c3",x"fe"),
   937 => (x"cd",x"02",x"99",x"49"),
   938 => (x"a9",x"ec",x"c0",x"87"),
   939 => (x"c0",x"87",x"c7",x"02"),
   940 => (x"ff",x"05",x"a9",x"fb"),
   941 => (x"66",x"d0",x"87",x"d5"),
   942 => (x"c0",x"87",x"c3",x"02"),
   943 => (x"ec",x"c0",x"7b",x"97"),
   944 => (x"87",x"c4",x"05",x"a9"),
   945 => (x"87",x"c5",x"4a",x"74"),
   946 => (x"0a",x"c0",x"4a",x"74"),
   947 => (x"c2",x"48",x"72",x"8a"),
   948 => (x"26",x"4d",x"26",x"87"),
   949 => (x"26",x"4b",x"26",x"4c"),
   950 => (x"c9",x"fd",x"1e",x"4f"),
   951 => (x"c0",x"49",x"70",x"87"),
   952 => (x"04",x"a9",x"b7",x"f0"),
   953 => (x"f9",x"c0",x"87",x"ca"),
   954 => (x"c3",x"01",x"a9",x"b7"),
   955 => (x"89",x"f0",x"c0",x"87"),
   956 => (x"a9",x"b7",x"c1",x"c1"),
   957 => (x"c1",x"87",x"ca",x"04"),
   958 => (x"01",x"a9",x"b7",x"da"),
   959 => (x"f7",x"c0",x"87",x"c3"),
   960 => (x"26",x"48",x"71",x"89"),
   961 => (x"5b",x"5e",x"0e",x"4f"),
   962 => (x"4a",x"71",x"0e",x"5c"),
   963 => (x"72",x"4c",x"d4",x"ff"),
   964 => (x"87",x"ea",x"c0",x"49"),
   965 => (x"02",x"9b",x"4b",x"70"),
   966 => (x"8b",x"c1",x"87",x"c2"),
   967 => (x"c8",x"48",x"d0",x"ff"),
   968 => (x"d5",x"c1",x"78",x"c5"),
   969 => (x"c6",x"49",x"73",x"7c"),
   970 => (x"fa",x"e0",x"c2",x"31"),
   971 => (x"48",x"4a",x"bf",x"97"),
   972 => (x"7c",x"70",x"b0",x"71"),
   973 => (x"c4",x"48",x"d0",x"ff"),
   974 => (x"fe",x"48",x"73",x"78"),
   975 => (x"5e",x"0e",x"87",x"d5"),
   976 => (x"0e",x"5d",x"5c",x"5b"),
   977 => (x"4c",x"71",x"86",x"f8"),
   978 => (x"e4",x"fb",x"7e",x"c0"),
   979 => (x"c0",x"4b",x"c0",x"87"),
   980 => (x"bf",x"97",x"eb",x"ff"),
   981 => (x"04",x"a9",x"c0",x"49"),
   982 => (x"f9",x"fb",x"87",x"cf"),
   983 => (x"c0",x"83",x"c1",x"87"),
   984 => (x"bf",x"97",x"eb",x"ff"),
   985 => (x"f1",x"06",x"ab",x"49"),
   986 => (x"eb",x"ff",x"c0",x"87"),
   987 => (x"cf",x"02",x"bf",x"97"),
   988 => (x"87",x"f2",x"fa",x"87"),
   989 => (x"02",x"99",x"49",x"70"),
   990 => (x"ec",x"c0",x"87",x"c6"),
   991 => (x"87",x"f1",x"05",x"a9"),
   992 => (x"e1",x"fa",x"4b",x"c0"),
   993 => (x"fa",x"4d",x"70",x"87"),
   994 => (x"a6",x"c8",x"87",x"dc"),
   995 => (x"87",x"d6",x"fa",x"58"),
   996 => (x"83",x"c1",x"4a",x"70"),
   997 => (x"97",x"49",x"a4",x"c8"),
   998 => (x"02",x"ad",x"49",x"69"),
   999 => (x"ff",x"c0",x"87",x"c7"),
  1000 => (x"e7",x"c0",x"05",x"ad"),
  1001 => (x"49",x"a4",x"c9",x"87"),
  1002 => (x"c4",x"49",x"69",x"97"),
  1003 => (x"c7",x"02",x"a9",x"66"),
  1004 => (x"ff",x"c0",x"48",x"87"),
  1005 => (x"87",x"d4",x"05",x"a8"),
  1006 => (x"97",x"49",x"a4",x"ca"),
  1007 => (x"02",x"aa",x"49",x"69"),
  1008 => (x"ff",x"c0",x"87",x"c6"),
  1009 => (x"87",x"c4",x"05",x"aa"),
  1010 => (x"87",x"d0",x"7e",x"c1"),
  1011 => (x"02",x"ad",x"ec",x"c0"),
  1012 => (x"fb",x"c0",x"87",x"c6"),
  1013 => (x"87",x"c4",x"05",x"ad"),
  1014 => (x"7e",x"c1",x"4b",x"c0"),
  1015 => (x"e1",x"fe",x"02",x"6e"),
  1016 => (x"87",x"e9",x"f9",x"87"),
  1017 => (x"8e",x"f8",x"48",x"73"),
  1018 => (x"00",x"87",x"e6",x"fb"),
  1019 => (x"5c",x"5b",x"5e",x"0e"),
  1020 => (x"71",x"1e",x"0e",x"5d"),
  1021 => (x"4d",x"4c",x"c0",x"4b"),
  1022 => (x"e8",x"c0",x"04",x"ab"),
  1023 => (x"fe",x"fc",x"c0",x"87"),
  1024 => (x"02",x"9d",x"75",x"1e"),
  1025 => (x"4a",x"c0",x"87",x"c4"),
  1026 => (x"4a",x"c1",x"87",x"c2"),
  1027 => (x"df",x"f0",x"49",x"72"),
  1028 => (x"70",x"86",x"c4",x"87"),
  1029 => (x"6e",x"84",x"c1",x"7e"),
  1030 => (x"73",x"87",x"c2",x"05"),
  1031 => (x"73",x"85",x"c1",x"4c"),
  1032 => (x"d8",x"ff",x"06",x"ac"),
  1033 => (x"26",x"48",x"6e",x"87"),
  1034 => (x"4c",x"26",x"4d",x"26"),
  1035 => (x"4f",x"26",x"4b",x"26"),
  1036 => (x"5c",x"5b",x"5e",x"0e"),
  1037 => (x"71",x"1e",x"0e",x"5d"),
  1038 => (x"91",x"de",x"49",x"4c"),
  1039 => (x"4d",x"c1",x"f0",x"c2"),
  1040 => (x"6d",x"97",x"85",x"71"),
  1041 => (x"87",x"dd",x"c1",x"02"),
  1042 => (x"bf",x"ec",x"ef",x"c2"),
  1043 => (x"72",x"82",x"74",x"4a"),
  1044 => (x"87",x"d8",x"fe",x"49"),
  1045 => (x"02",x"6e",x"7e",x"70"),
  1046 => (x"c2",x"87",x"f3",x"c0"),
  1047 => (x"6e",x"4b",x"f4",x"ef"),
  1048 => (x"ff",x"49",x"cb",x"4a"),
  1049 => (x"74",x"87",x"c1",x"c1"),
  1050 => (x"c1",x"93",x"cb",x"4b"),
  1051 => (x"c4",x"83",x"dd",x"e3"),
  1052 => (x"e9",x"c2",x"c1",x"83"),
  1053 => (x"c1",x"49",x"74",x"7b"),
  1054 => (x"75",x"87",x"d1",x"c3"),
  1055 => (x"c0",x"f0",x"c2",x"7b"),
  1056 => (x"1e",x"49",x"bf",x"97"),
  1057 => (x"49",x"f4",x"ef",x"c2"),
  1058 => (x"87",x"f0",x"dd",x"c1"),
  1059 => (x"49",x"74",x"86",x"c4"),
  1060 => (x"87",x"f8",x"c2",x"c1"),
  1061 => (x"c4",x"c1",x"49",x"c0"),
  1062 => (x"ef",x"c2",x"87",x"d7"),
  1063 => (x"78",x"c0",x"48",x"e8"),
  1064 => (x"cb",x"dd",x"49",x"c1"),
  1065 => (x"ff",x"fd",x"26",x"87"),
  1066 => (x"61",x"6f",x"4c",x"87"),
  1067 => (x"67",x"6e",x"69",x"64"),
  1068 => (x"00",x"2e",x"2e",x"2e"),
  1069 => (x"5c",x"5b",x"5e",x"0e"),
  1070 => (x"4a",x"4b",x"71",x"0e"),
  1071 => (x"bf",x"ec",x"ef",x"c2"),
  1072 => (x"fc",x"49",x"72",x"82"),
  1073 => (x"4c",x"70",x"87",x"e6"),
  1074 => (x"87",x"c4",x"02",x"9c"),
  1075 => (x"87",x"e8",x"ec",x"49"),
  1076 => (x"48",x"ec",x"ef",x"c2"),
  1077 => (x"49",x"c1",x"78",x"c0"),
  1078 => (x"fd",x"87",x"d5",x"dc"),
  1079 => (x"5e",x"0e",x"87",x"cc"),
  1080 => (x"0e",x"5d",x"5c",x"5b"),
  1081 => (x"e2",x"c2",x"86",x"f4"),
  1082 => (x"4c",x"c0",x"4d",x"f6"),
  1083 => (x"c0",x"48",x"a6",x"c4"),
  1084 => (x"ec",x"ef",x"c2",x"78"),
  1085 => (x"a9",x"c0",x"49",x"bf"),
  1086 => (x"87",x"c1",x"c1",x"06"),
  1087 => (x"48",x"f6",x"e2",x"c2"),
  1088 => (x"f8",x"c0",x"02",x"98"),
  1089 => (x"fe",x"fc",x"c0",x"87"),
  1090 => (x"02",x"66",x"c8",x"1e"),
  1091 => (x"a6",x"c4",x"87",x"c7"),
  1092 => (x"c5",x"78",x"c0",x"48"),
  1093 => (x"48",x"a6",x"c4",x"87"),
  1094 => (x"66",x"c4",x"78",x"c1"),
  1095 => (x"87",x"d0",x"ec",x"49"),
  1096 => (x"4d",x"70",x"86",x"c4"),
  1097 => (x"66",x"c4",x"84",x"c1"),
  1098 => (x"c8",x"80",x"c1",x"48"),
  1099 => (x"ef",x"c2",x"58",x"a6"),
  1100 => (x"ac",x"49",x"bf",x"ec"),
  1101 => (x"75",x"87",x"c6",x"03"),
  1102 => (x"c8",x"ff",x"05",x"9d"),
  1103 => (x"75",x"4c",x"c0",x"87"),
  1104 => (x"e0",x"c3",x"02",x"9d"),
  1105 => (x"fe",x"fc",x"c0",x"87"),
  1106 => (x"02",x"66",x"c8",x"1e"),
  1107 => (x"a6",x"cc",x"87",x"c7"),
  1108 => (x"c5",x"78",x"c0",x"48"),
  1109 => (x"48",x"a6",x"cc",x"87"),
  1110 => (x"66",x"cc",x"78",x"c1"),
  1111 => (x"87",x"d0",x"eb",x"49"),
  1112 => (x"7e",x"70",x"86",x"c4"),
  1113 => (x"e9",x"c2",x"02",x"6e"),
  1114 => (x"cb",x"49",x"6e",x"87"),
  1115 => (x"49",x"69",x"97",x"81"),
  1116 => (x"c1",x"02",x"99",x"d0"),
  1117 => (x"c2",x"c1",x"87",x"d6"),
  1118 => (x"49",x"74",x"4a",x"f4"),
  1119 => (x"e3",x"c1",x"91",x"cb"),
  1120 => (x"79",x"72",x"81",x"dd"),
  1121 => (x"ff",x"c3",x"81",x"c8"),
  1122 => (x"de",x"49",x"74",x"51"),
  1123 => (x"c1",x"f0",x"c2",x"91"),
  1124 => (x"c2",x"85",x"71",x"4d"),
  1125 => (x"c1",x"7d",x"97",x"c1"),
  1126 => (x"e0",x"c0",x"49",x"a5"),
  1127 => (x"c6",x"eb",x"c2",x"51"),
  1128 => (x"d2",x"02",x"bf",x"97"),
  1129 => (x"c2",x"84",x"c1",x"87"),
  1130 => (x"eb",x"c2",x"4b",x"a5"),
  1131 => (x"49",x"db",x"4a",x"c6"),
  1132 => (x"87",x"f4",x"fb",x"fe"),
  1133 => (x"cd",x"87",x"db",x"c1"),
  1134 => (x"51",x"c0",x"49",x"a5"),
  1135 => (x"a5",x"c2",x"84",x"c1"),
  1136 => (x"cb",x"4a",x"6e",x"4b"),
  1137 => (x"df",x"fb",x"fe",x"49"),
  1138 => (x"87",x"c6",x"c1",x"87"),
  1139 => (x"4a",x"f0",x"c0",x"c1"),
  1140 => (x"91",x"cb",x"49",x"74"),
  1141 => (x"81",x"dd",x"e3",x"c1"),
  1142 => (x"eb",x"c2",x"79",x"72"),
  1143 => (x"02",x"bf",x"97",x"c6"),
  1144 => (x"49",x"74",x"87",x"d8"),
  1145 => (x"84",x"c1",x"91",x"de"),
  1146 => (x"4b",x"c1",x"f0",x"c2"),
  1147 => (x"eb",x"c2",x"83",x"71"),
  1148 => (x"49",x"dd",x"4a",x"c6"),
  1149 => (x"87",x"f0",x"fa",x"fe"),
  1150 => (x"4b",x"74",x"87",x"d8"),
  1151 => (x"f0",x"c2",x"93",x"de"),
  1152 => (x"a3",x"cb",x"83",x"c1"),
  1153 => (x"c1",x"51",x"c0",x"49"),
  1154 => (x"4a",x"6e",x"73",x"84"),
  1155 => (x"fa",x"fe",x"49",x"cb"),
  1156 => (x"66",x"c4",x"87",x"d6"),
  1157 => (x"c8",x"80",x"c1",x"48"),
  1158 => (x"ac",x"c7",x"58",x"a6"),
  1159 => (x"87",x"c5",x"c0",x"03"),
  1160 => (x"e0",x"fc",x"05",x"6e"),
  1161 => (x"f4",x"48",x"74",x"87"),
  1162 => (x"87",x"fc",x"f7",x"8e"),
  1163 => (x"71",x"1e",x"73",x"1e"),
  1164 => (x"91",x"cb",x"49",x"4b"),
  1165 => (x"81",x"dd",x"e3",x"c1"),
  1166 => (x"c2",x"4a",x"a1",x"c8"),
  1167 => (x"12",x"48",x"fa",x"e0"),
  1168 => (x"4a",x"a1",x"c9",x"50"),
  1169 => (x"48",x"eb",x"ff",x"c0"),
  1170 => (x"81",x"ca",x"50",x"12"),
  1171 => (x"48",x"c0",x"f0",x"c2"),
  1172 => (x"f0",x"c2",x"50",x"11"),
  1173 => (x"49",x"bf",x"97",x"c0"),
  1174 => (x"c1",x"49",x"c0",x"1e"),
  1175 => (x"c2",x"87",x"dd",x"d6"),
  1176 => (x"de",x"48",x"e8",x"ef"),
  1177 => (x"d6",x"49",x"c1",x"78"),
  1178 => (x"f6",x"26",x"87",x"c6"),
  1179 => (x"71",x"1e",x"87",x"fe"),
  1180 => (x"91",x"cb",x"49",x"4a"),
  1181 => (x"81",x"dd",x"e3",x"c1"),
  1182 => (x"48",x"11",x"81",x"c8"),
  1183 => (x"58",x"ec",x"ef",x"c2"),
  1184 => (x"48",x"ec",x"ef",x"c2"),
  1185 => (x"49",x"c1",x"78",x"c0"),
  1186 => (x"26",x"87",x"e5",x"d5"),
  1187 => (x"49",x"c0",x"1e",x"4f"),
  1188 => (x"87",x"dd",x"fc",x"c0"),
  1189 => (x"71",x"1e",x"4f",x"26"),
  1190 => (x"87",x"d2",x"02",x"99"),
  1191 => (x"48",x"f2",x"e4",x"c1"),
  1192 => (x"80",x"f7",x"50",x"c0"),
  1193 => (x"40",x"ee",x"c9",x"c1"),
  1194 => (x"78",x"d6",x"e3",x"c1"),
  1195 => (x"e4",x"c1",x"87",x"ce"),
  1196 => (x"e3",x"c1",x"48",x"ee"),
  1197 => (x"80",x"fc",x"78",x"cf"),
  1198 => (x"78",x"cd",x"ca",x"c1"),
  1199 => (x"5e",x"0e",x"4f",x"26"),
  1200 => (x"71",x"0e",x"5c",x"5b"),
  1201 => (x"92",x"cb",x"4a",x"4c"),
  1202 => (x"82",x"dd",x"e3",x"c1"),
  1203 => (x"c9",x"49",x"a2",x"c8"),
  1204 => (x"6b",x"97",x"4b",x"a2"),
  1205 => (x"69",x"97",x"1e",x"4b"),
  1206 => (x"82",x"ca",x"1e",x"49"),
  1207 => (x"e7",x"c0",x"49",x"12"),
  1208 => (x"49",x"c0",x"87",x"d8"),
  1209 => (x"74",x"87",x"c9",x"d4"),
  1210 => (x"df",x"f9",x"c0",x"49"),
  1211 => (x"f4",x"8e",x"f8",x"87"),
  1212 => (x"73",x"1e",x"87",x"f8"),
  1213 => (x"49",x"4b",x"71",x"1e"),
  1214 => (x"73",x"87",x"c3",x"ff"),
  1215 => (x"87",x"fe",x"fe",x"49"),
  1216 => (x"1e",x"87",x"e9",x"f4"),
  1217 => (x"4b",x"71",x"1e",x"73"),
  1218 => (x"02",x"4a",x"a3",x"c6"),
  1219 => (x"8a",x"c1",x"87",x"db"),
  1220 => (x"8a",x"87",x"d6",x"02"),
  1221 => (x"87",x"da",x"c1",x"02"),
  1222 => (x"fc",x"c0",x"02",x"8a"),
  1223 => (x"c0",x"02",x"8a",x"87"),
  1224 => (x"02",x"8a",x"87",x"e1"),
  1225 => (x"db",x"c1",x"87",x"cb"),
  1226 => (x"fd",x"49",x"c7",x"87"),
  1227 => (x"de",x"c1",x"87",x"c0"),
  1228 => (x"ec",x"ef",x"c2",x"87"),
  1229 => (x"cb",x"c1",x"02",x"bf"),
  1230 => (x"88",x"c1",x"48",x"87"),
  1231 => (x"58",x"f0",x"ef",x"c2"),
  1232 => (x"c2",x"87",x"c1",x"c1"),
  1233 => (x"02",x"bf",x"f0",x"ef"),
  1234 => (x"c2",x"87",x"f9",x"c0"),
  1235 => (x"48",x"bf",x"ec",x"ef"),
  1236 => (x"ef",x"c2",x"80",x"c1"),
  1237 => (x"eb",x"c0",x"58",x"f0"),
  1238 => (x"ec",x"ef",x"c2",x"87"),
  1239 => (x"89",x"c6",x"49",x"bf"),
  1240 => (x"59",x"f0",x"ef",x"c2"),
  1241 => (x"03",x"a9",x"b7",x"c0"),
  1242 => (x"ef",x"c2",x"87",x"da"),
  1243 => (x"78",x"c0",x"48",x"ec"),
  1244 => (x"ef",x"c2",x"87",x"d2"),
  1245 => (x"cb",x"02",x"bf",x"f0"),
  1246 => (x"ec",x"ef",x"c2",x"87"),
  1247 => (x"80",x"c6",x"48",x"bf"),
  1248 => (x"58",x"f0",x"ef",x"c2"),
  1249 => (x"e7",x"d1",x"49",x"c0"),
  1250 => (x"c0",x"49",x"73",x"87"),
  1251 => (x"f2",x"87",x"fd",x"f6"),
  1252 => (x"5e",x"0e",x"87",x"da"),
  1253 => (x"71",x"0e",x"5c",x"5b"),
  1254 => (x"1e",x"66",x"cc",x"4c"),
  1255 => (x"93",x"cb",x"4b",x"74"),
  1256 => (x"83",x"dd",x"e3",x"c1"),
  1257 => (x"6a",x"4a",x"a3",x"c4"),
  1258 => (x"cb",x"f4",x"fe",x"49"),
  1259 => (x"ec",x"c8",x"c1",x"87"),
  1260 => (x"49",x"a3",x"c8",x"7b"),
  1261 => (x"c9",x"51",x"66",x"d4"),
  1262 => (x"66",x"d8",x"49",x"a3"),
  1263 => (x"49",x"a3",x"ca",x"51"),
  1264 => (x"26",x"51",x"66",x"dc"),
  1265 => (x"0e",x"87",x"e3",x"f1"),
  1266 => (x"5d",x"5c",x"5b",x"5e"),
  1267 => (x"86",x"d0",x"ff",x"0e"),
  1268 => (x"c4",x"59",x"a6",x"d8"),
  1269 => (x"78",x"c0",x"48",x"a6"),
  1270 => (x"c4",x"c1",x"80",x"c4"),
  1271 => (x"80",x"c4",x"78",x"66"),
  1272 => (x"80",x"c4",x"78",x"c1"),
  1273 => (x"ef",x"c2",x"78",x"c1"),
  1274 => (x"78",x"c1",x"48",x"f0"),
  1275 => (x"bf",x"e8",x"ef",x"c2"),
  1276 => (x"05",x"a8",x"de",x"48"),
  1277 => (x"e5",x"f3",x"87",x"cb"),
  1278 => (x"c8",x"49",x"70",x"87"),
  1279 => (x"f8",x"ce",x"59",x"a6"),
  1280 => (x"87",x"ed",x"e8",x"87"),
  1281 => (x"e8",x"87",x"cf",x"e9"),
  1282 => (x"4c",x"70",x"87",x"dc"),
  1283 => (x"02",x"ac",x"fb",x"c0"),
  1284 => (x"d4",x"87",x"d0",x"c1"),
  1285 => (x"c2",x"c1",x"05",x"66"),
  1286 => (x"1e",x"1e",x"c0",x"87"),
  1287 => (x"e5",x"c1",x"1e",x"c1"),
  1288 => (x"49",x"c0",x"1e",x"d0"),
  1289 => (x"c1",x"87",x"eb",x"fd"),
  1290 => (x"c4",x"4a",x"66",x"d0"),
  1291 => (x"c7",x"49",x"6a",x"82"),
  1292 => (x"c1",x"51",x"74",x"81"),
  1293 => (x"6a",x"1e",x"d8",x"1e"),
  1294 => (x"e8",x"81",x"c8",x"49"),
  1295 => (x"86",x"d8",x"87",x"ec"),
  1296 => (x"48",x"66",x"c4",x"c1"),
  1297 => (x"c7",x"01",x"a8",x"c0"),
  1298 => (x"48",x"a6",x"c4",x"87"),
  1299 => (x"87",x"ce",x"78",x"c1"),
  1300 => (x"48",x"66",x"c4",x"c1"),
  1301 => (x"a6",x"cc",x"88",x"c1"),
  1302 => (x"e7",x"87",x"c3",x"58"),
  1303 => (x"a6",x"cc",x"87",x"f8"),
  1304 => (x"74",x"78",x"c2",x"48"),
  1305 => (x"cc",x"cd",x"02",x"9c"),
  1306 => (x"48",x"66",x"c4",x"87"),
  1307 => (x"a8",x"66",x"c8",x"c1"),
  1308 => (x"87",x"c1",x"cd",x"03"),
  1309 => (x"c0",x"48",x"a6",x"d8"),
  1310 => (x"87",x"ea",x"e6",x"78"),
  1311 => (x"d0",x"c1",x"4c",x"70"),
  1312 => (x"d6",x"c2",x"05",x"ac"),
  1313 => (x"7e",x"66",x"d8",x"87"),
  1314 => (x"70",x"87",x"ce",x"e9"),
  1315 => (x"59",x"a6",x"dc",x"49"),
  1316 => (x"70",x"87",x"d3",x"e6"),
  1317 => (x"ac",x"ec",x"c0",x"4c"),
  1318 => (x"87",x"ea",x"c1",x"05"),
  1319 => (x"cb",x"49",x"66",x"c4"),
  1320 => (x"66",x"c0",x"c1",x"91"),
  1321 => (x"4a",x"a1",x"c4",x"81"),
  1322 => (x"a1",x"c8",x"4d",x"6a"),
  1323 => (x"52",x"66",x"d8",x"4a"),
  1324 => (x"79",x"ee",x"c9",x"c1"),
  1325 => (x"70",x"87",x"ef",x"e5"),
  1326 => (x"d8",x"02",x"9c",x"4c"),
  1327 => (x"ac",x"fb",x"c0",x"87"),
  1328 => (x"74",x"87",x"d2",x"02"),
  1329 => (x"87",x"de",x"e5",x"55"),
  1330 => (x"02",x"9c",x"4c",x"70"),
  1331 => (x"fb",x"c0",x"87",x"c7"),
  1332 => (x"ee",x"ff",x"05",x"ac"),
  1333 => (x"55",x"e0",x"c0",x"87"),
  1334 => (x"c0",x"55",x"c1",x"c2"),
  1335 => (x"66",x"d4",x"7d",x"97"),
  1336 => (x"05",x"a9",x"6e",x"49"),
  1337 => (x"66",x"c4",x"87",x"db"),
  1338 => (x"a8",x"66",x"c8",x"48"),
  1339 => (x"c4",x"87",x"ca",x"04"),
  1340 => (x"80",x"c1",x"48",x"66"),
  1341 => (x"c8",x"58",x"a6",x"c8"),
  1342 => (x"48",x"66",x"c8",x"87"),
  1343 => (x"a6",x"cc",x"88",x"c1"),
  1344 => (x"87",x"e2",x"e4",x"58"),
  1345 => (x"d0",x"c1",x"4c",x"70"),
  1346 => (x"87",x"c8",x"05",x"ac"),
  1347 => (x"c1",x"48",x"66",x"d0"),
  1348 => (x"58",x"a6",x"d4",x"80"),
  1349 => (x"02",x"ac",x"d0",x"c1"),
  1350 => (x"dc",x"87",x"ea",x"fd"),
  1351 => (x"66",x"d4",x"48",x"a6"),
  1352 => (x"48",x"66",x"d8",x"78"),
  1353 => (x"05",x"a8",x"66",x"dc"),
  1354 => (x"c0",x"87",x"dc",x"c9"),
  1355 => (x"c0",x"48",x"a6",x"e0"),
  1356 => (x"80",x"c4",x"78",x"f0"),
  1357 => (x"c4",x"78",x"66",x"cc"),
  1358 => (x"7e",x"78",x"c0",x"80"),
  1359 => (x"fb",x"c0",x"48",x"74"),
  1360 => (x"a6",x"f0",x"c0",x"88"),
  1361 => (x"02",x"98",x"70",x"58"),
  1362 => (x"48",x"87",x"d7",x"c8"),
  1363 => (x"f0",x"c0",x"88",x"cb"),
  1364 => (x"98",x"70",x"58",x"a6"),
  1365 => (x"87",x"e9",x"c0",x"02"),
  1366 => (x"c0",x"88",x"c9",x"48"),
  1367 => (x"70",x"58",x"a6",x"f0"),
  1368 => (x"e1",x"c3",x"02",x"98"),
  1369 => (x"88",x"c4",x"48",x"87"),
  1370 => (x"58",x"a6",x"f0",x"c0"),
  1371 => (x"de",x"02",x"98",x"70"),
  1372 => (x"88",x"c1",x"48",x"87"),
  1373 => (x"58",x"a6",x"f0",x"c0"),
  1374 => (x"c3",x"02",x"98",x"70"),
  1375 => (x"db",x"c7",x"87",x"c8"),
  1376 => (x"a6",x"e0",x"c0",x"87"),
  1377 => (x"cc",x"78",x"c0",x"48"),
  1378 => (x"80",x"c1",x"48",x"66"),
  1379 => (x"e2",x"58",x"a6",x"d0"),
  1380 => (x"4c",x"70",x"87",x"d4"),
  1381 => (x"02",x"ac",x"ec",x"c0"),
  1382 => (x"e0",x"c0",x"87",x"d5"),
  1383 => (x"87",x"c6",x"02",x"66"),
  1384 => (x"5c",x"a6",x"e4",x"c0"),
  1385 => (x"48",x"74",x"87",x"c9"),
  1386 => (x"c0",x"88",x"f0",x"c0"),
  1387 => (x"c0",x"58",x"a6",x"e8"),
  1388 => (x"cc",x"02",x"ac",x"ec"),
  1389 => (x"87",x"ee",x"e1",x"87"),
  1390 => (x"ec",x"c0",x"4c",x"70"),
  1391 => (x"f4",x"ff",x"05",x"ac"),
  1392 => (x"66",x"e0",x"c0",x"87"),
  1393 => (x"49",x"66",x"d4",x"1e"),
  1394 => (x"66",x"ec",x"c0",x"1e"),
  1395 => (x"d0",x"e5",x"c1",x"1e"),
  1396 => (x"49",x"66",x"d4",x"1e"),
  1397 => (x"c0",x"87",x"fb",x"f6"),
  1398 => (x"dc",x"1e",x"ca",x"1e"),
  1399 => (x"91",x"cb",x"49",x"66"),
  1400 => (x"81",x"66",x"d8",x"c1"),
  1401 => (x"c4",x"48",x"a6",x"d8"),
  1402 => (x"66",x"d8",x"78",x"a1"),
  1403 => (x"f9",x"e1",x"49",x"bf"),
  1404 => (x"c0",x"86",x"d8",x"87"),
  1405 => (x"c1",x"06",x"a8",x"b7"),
  1406 => (x"1e",x"c1",x"87",x"c7"),
  1407 => (x"66",x"c8",x"1e",x"de"),
  1408 => (x"e5",x"e1",x"49",x"bf"),
  1409 => (x"70",x"86",x"c8",x"87"),
  1410 => (x"08",x"c0",x"48",x"49"),
  1411 => (x"a6",x"e4",x"c0",x"88"),
  1412 => (x"a8",x"b7",x"c0",x"58"),
  1413 => (x"87",x"e9",x"c0",x"06"),
  1414 => (x"48",x"66",x"e0",x"c0"),
  1415 => (x"03",x"a8",x"b7",x"dd"),
  1416 => (x"bf",x"6e",x"87",x"df"),
  1417 => (x"66",x"e0",x"c0",x"49"),
  1418 => (x"51",x"e0",x"c0",x"81"),
  1419 => (x"81",x"c1",x"49",x"66"),
  1420 => (x"c2",x"81",x"bf",x"6e"),
  1421 => (x"e0",x"c0",x"51",x"c1"),
  1422 => (x"81",x"c2",x"49",x"66"),
  1423 => (x"c0",x"81",x"bf",x"6e"),
  1424 => (x"c4",x"7e",x"c1",x"51"),
  1425 => (x"d0",x"e2",x"87",x"dc"),
  1426 => (x"a6",x"e4",x"c0",x"87"),
  1427 => (x"87",x"c9",x"e2",x"58"),
  1428 => (x"58",x"a6",x"e8",x"c0"),
  1429 => (x"05",x"a8",x"ec",x"c0"),
  1430 => (x"c0",x"87",x"cb",x"c0"),
  1431 => (x"c0",x"48",x"a6",x"e4"),
  1432 => (x"c0",x"78",x"66",x"e0"),
  1433 => (x"de",x"ff",x"87",x"c4"),
  1434 => (x"66",x"c4",x"87",x"fc"),
  1435 => (x"c1",x"91",x"cb",x"49"),
  1436 => (x"71",x"48",x"66",x"c0"),
  1437 => (x"6e",x"7e",x"70",x"80"),
  1438 => (x"6e",x"82",x"c8",x"4a"),
  1439 => (x"c0",x"81",x"ca",x"49"),
  1440 => (x"c0",x"51",x"66",x"e0"),
  1441 => (x"c1",x"49",x"66",x"e4"),
  1442 => (x"66",x"e0",x"c0",x"81"),
  1443 => (x"71",x"48",x"c1",x"89"),
  1444 => (x"c1",x"49",x"70",x"30"),
  1445 => (x"7a",x"97",x"71",x"89"),
  1446 => (x"bf",x"dd",x"f3",x"c2"),
  1447 => (x"66",x"e0",x"c0",x"49"),
  1448 => (x"4a",x"6a",x"97",x"29"),
  1449 => (x"c0",x"98",x"71",x"48"),
  1450 => (x"6e",x"58",x"a6",x"f0"),
  1451 => (x"69",x"81",x"c4",x"49"),
  1452 => (x"48",x"66",x"dc",x"4d"),
  1453 => (x"02",x"a8",x"66",x"d8"),
  1454 => (x"d8",x"87",x"c8",x"c0"),
  1455 => (x"78",x"c0",x"48",x"a6"),
  1456 => (x"d8",x"87",x"c5",x"c0"),
  1457 => (x"78",x"c1",x"48",x"a6"),
  1458 => (x"c0",x"1e",x"66",x"d8"),
  1459 => (x"49",x"75",x"1e",x"e0"),
  1460 => (x"87",x"d6",x"de",x"ff"),
  1461 => (x"4c",x"70",x"86",x"c8"),
  1462 => (x"06",x"ac",x"b7",x"c0"),
  1463 => (x"74",x"87",x"d4",x"c1"),
  1464 => (x"49",x"e0",x"c0",x"85"),
  1465 => (x"4b",x"75",x"89",x"74"),
  1466 => (x"4a",x"ed",x"df",x"c1"),
  1467 => (x"f7",x"e6",x"fe",x"71"),
  1468 => (x"c0",x"85",x"c2",x"87"),
  1469 => (x"c1",x"48",x"66",x"e8"),
  1470 => (x"a6",x"ec",x"c0",x"80"),
  1471 => (x"66",x"ec",x"c0",x"58"),
  1472 => (x"70",x"81",x"c1",x"49"),
  1473 => (x"c8",x"c0",x"02",x"a9"),
  1474 => (x"48",x"a6",x"d8",x"87"),
  1475 => (x"c5",x"c0",x"78",x"c0"),
  1476 => (x"48",x"a6",x"d8",x"87"),
  1477 => (x"66",x"d8",x"78",x"c1"),
  1478 => (x"49",x"a4",x"c2",x"1e"),
  1479 => (x"71",x"48",x"e0",x"c0"),
  1480 => (x"1e",x"49",x"70",x"88"),
  1481 => (x"dd",x"ff",x"49",x"75"),
  1482 => (x"86",x"c8",x"87",x"c0"),
  1483 => (x"01",x"a8",x"b7",x"c0"),
  1484 => (x"c0",x"87",x"c0",x"ff"),
  1485 => (x"c0",x"02",x"66",x"e8"),
  1486 => (x"49",x"6e",x"87",x"d1"),
  1487 => (x"e8",x"c0",x"81",x"c9"),
  1488 => (x"48",x"6e",x"51",x"66"),
  1489 => (x"78",x"fe",x"ca",x"c1"),
  1490 => (x"6e",x"87",x"cc",x"c0"),
  1491 => (x"c2",x"81",x"c9",x"49"),
  1492 => (x"c1",x"48",x"6e",x"51"),
  1493 => (x"c1",x"78",x"f2",x"cb"),
  1494 => (x"87",x"c6",x"c0",x"7e"),
  1495 => (x"87",x"f6",x"db",x"ff"),
  1496 => (x"02",x"6e",x"4c",x"70"),
  1497 => (x"c4",x"87",x"f5",x"c0"),
  1498 => (x"66",x"c8",x"48",x"66"),
  1499 => (x"cb",x"c0",x"04",x"a8"),
  1500 => (x"48",x"66",x"c4",x"87"),
  1501 => (x"a6",x"c8",x"80",x"c1"),
  1502 => (x"87",x"e0",x"c0",x"58"),
  1503 => (x"c1",x"48",x"66",x"c8"),
  1504 => (x"58",x"a6",x"cc",x"88"),
  1505 => (x"c1",x"87",x"d5",x"c0"),
  1506 => (x"c0",x"05",x"ac",x"c6"),
  1507 => (x"66",x"cc",x"87",x"c8"),
  1508 => (x"d0",x"80",x"c1",x"48"),
  1509 => (x"da",x"ff",x"58",x"a6"),
  1510 => (x"4c",x"70",x"87",x"fc"),
  1511 => (x"c1",x"48",x"66",x"d0"),
  1512 => (x"58",x"a6",x"d4",x"80"),
  1513 => (x"c0",x"02",x"9c",x"74"),
  1514 => (x"66",x"c4",x"87",x"cb"),
  1515 => (x"66",x"c8",x"c1",x"48"),
  1516 => (x"ff",x"f2",x"04",x"a8"),
  1517 => (x"d4",x"da",x"ff",x"87"),
  1518 => (x"48",x"66",x"c4",x"87"),
  1519 => (x"c0",x"03",x"a8",x"c7"),
  1520 => (x"ef",x"c2",x"87",x"e5"),
  1521 => (x"78",x"c0",x"48",x"f0"),
  1522 => (x"cb",x"49",x"66",x"c4"),
  1523 => (x"66",x"c0",x"c1",x"91"),
  1524 => (x"4a",x"a1",x"c4",x"81"),
  1525 => (x"52",x"c0",x"4a",x"6a"),
  1526 => (x"48",x"66",x"c4",x"79"),
  1527 => (x"a6",x"c8",x"80",x"c1"),
  1528 => (x"04",x"a8",x"c7",x"58"),
  1529 => (x"ff",x"87",x"db",x"ff"),
  1530 => (x"fb",x"e0",x"8e",x"d0"),
  1531 => (x"00",x"20",x"3a",x"87"),
  1532 => (x"71",x"1e",x"73",x"1e"),
  1533 => (x"c6",x"02",x"9b",x"4b"),
  1534 => (x"ec",x"ef",x"c2",x"87"),
  1535 => (x"c7",x"78",x"c0",x"48"),
  1536 => (x"ec",x"ef",x"c2",x"1e"),
  1537 => (x"c1",x"1e",x"49",x"bf"),
  1538 => (x"c2",x"1e",x"dd",x"e3"),
  1539 => (x"49",x"bf",x"e8",x"ef"),
  1540 => (x"cc",x"87",x"f4",x"ee"),
  1541 => (x"e8",x"ef",x"c2",x"86"),
  1542 => (x"f9",x"e9",x"49",x"bf"),
  1543 => (x"02",x"9b",x"73",x"87"),
  1544 => (x"e3",x"c1",x"87",x"c8"),
  1545 => (x"e5",x"c0",x"49",x"dd"),
  1546 => (x"df",x"ff",x"87",x"f4"),
  1547 => (x"c2",x"1e",x"87",x"fe"),
  1548 => (x"c0",x"48",x"fa",x"e0"),
  1549 => (x"c0",x"e5",x"c1",x"50"),
  1550 => (x"fb",x"c0",x"49",x"bf"),
  1551 => (x"48",x"c0",x"87",x"d1"),
  1552 => (x"c7",x"1e",x"4f",x"26"),
  1553 => (x"49",x"c1",x"87",x"e9"),
  1554 => (x"fe",x"87",x"e5",x"fe"),
  1555 => (x"70",x"87",x"ec",x"e9"),
  1556 => (x"87",x"cd",x"02",x"98"),
  1557 => (x"87",x"e9",x"f2",x"fe"),
  1558 => (x"c4",x"02",x"98",x"70"),
  1559 => (x"c2",x"4a",x"c1",x"87"),
  1560 => (x"72",x"4a",x"c0",x"87"),
  1561 => (x"87",x"ce",x"05",x"9a"),
  1562 => (x"e2",x"c1",x"1e",x"c0"),
  1563 => (x"f0",x"c0",x"49",x"d6"),
  1564 => (x"86",x"c4",x"87",x"fb"),
  1565 => (x"ff",x"c0",x"87",x"fe"),
  1566 => (x"1e",x"c0",x"87",x"ea"),
  1567 => (x"49",x"e1",x"e2",x"c1"),
  1568 => (x"87",x"e9",x"f0",x"c0"),
  1569 => (x"e5",x"fe",x"1e",x"c0"),
  1570 => (x"c0",x"49",x"70",x"87"),
  1571 => (x"c3",x"87",x"de",x"f0"),
  1572 => (x"8e",x"f8",x"87",x"dc"),
  1573 => (x"44",x"53",x"4f",x"26"),
  1574 => (x"69",x"61",x"66",x"20"),
  1575 => (x"2e",x"64",x"65",x"6c"),
  1576 => (x"6f",x"6f",x"42",x"00"),
  1577 => (x"67",x"6e",x"69",x"74"),
  1578 => (x"00",x"2e",x"2e",x"2e"),
  1579 => (x"c9",x"e8",x"c0",x"1e"),
  1580 => (x"ee",x"f3",x"c0",x"87"),
  1581 => (x"26",x"87",x"f6",x"87"),
  1582 => (x"ef",x"c2",x"1e",x"4f"),
  1583 => (x"78",x"c0",x"48",x"ec"),
  1584 => (x"48",x"e8",x"ef",x"c2"),
  1585 => (x"f9",x"fd",x"78",x"c0"),
  1586 => (x"c0",x"87",x"e1",x"87"),
  1587 => (x"80",x"4f",x"26",x"48"),
  1588 => (x"69",x"78",x"45",x"20"),
  1589 => (x"20",x"80",x"00",x"74"),
  1590 => (x"6b",x"63",x"61",x"42"),
  1591 => (x"00",x"12",x"6e",x"00"),
  1592 => (x"00",x"2c",x"01",x"00"),
  1593 => (x"00",x"00",x"00",x"00"),
  1594 => (x"00",x"00",x"12",x"6e"),
  1595 => (x"00",x"00",x"2c",x"1f"),
  1596 => (x"6e",x"00",x"00",x"00"),
  1597 => (x"3d",x"00",x"00",x"12"),
  1598 => (x"00",x"00",x"00",x"2c"),
  1599 => (x"12",x"6e",x"00",x"00"),
  1600 => (x"2c",x"5b",x"00",x"00"),
  1601 => (x"00",x"00",x"00",x"00"),
  1602 => (x"00",x"12",x"6e",x"00"),
  1603 => (x"00",x"2c",x"79",x"00"),
  1604 => (x"00",x"00",x"00",x"00"),
  1605 => (x"00",x"00",x"12",x"6e"),
  1606 => (x"00",x"00",x"2c",x"97"),
  1607 => (x"6e",x"00",x"00",x"00"),
  1608 => (x"b5",x"00",x"00",x"12"),
  1609 => (x"00",x"00",x"00",x"2c"),
  1610 => (x"12",x"6e",x"00",x"00"),
  1611 => (x"00",x"00",x"00",x"00"),
  1612 => (x"00",x"00",x"00",x"00"),
  1613 => (x"00",x"13",x"03",x"00"),
  1614 => (x"00",x"00",x"00",x"00"),
  1615 => (x"00",x"00",x"00",x"00"),
  1616 => (x"00",x"00",x"19",x"44"),
  1617 => (x"54",x"4f",x"4f",x"42"),
  1618 => (x"20",x"20",x"20",x"20"),
  1619 => (x"00",x"4d",x"4f",x"52"),
  1620 => (x"64",x"61",x"6f",x"4c"),
  1621 => (x"00",x"2e",x"2a",x"20"),
  1622 => (x"48",x"f0",x"fe",x"1e"),
  1623 => (x"09",x"cd",x"78",x"c0"),
  1624 => (x"4f",x"26",x"09",x"79"),
  1625 => (x"f0",x"fe",x"1e",x"1e"),
  1626 => (x"26",x"48",x"7e",x"bf"),
  1627 => (x"fe",x"1e",x"4f",x"26"),
  1628 => (x"78",x"c1",x"48",x"f0"),
  1629 => (x"fe",x"1e",x"4f",x"26"),
  1630 => (x"78",x"c0",x"48",x"f0"),
  1631 => (x"71",x"1e",x"4f",x"26"),
  1632 => (x"52",x"52",x"c0",x"4a"),
  1633 => (x"5e",x"0e",x"4f",x"26"),
  1634 => (x"0e",x"5d",x"5c",x"5b"),
  1635 => (x"4d",x"71",x"86",x"f4"),
  1636 => (x"c1",x"7e",x"6d",x"97"),
  1637 => (x"6c",x"97",x"4c",x"a5"),
  1638 => (x"58",x"a6",x"c8",x"48"),
  1639 => (x"66",x"c4",x"48",x"6e"),
  1640 => (x"87",x"c5",x"05",x"a8"),
  1641 => (x"e6",x"c0",x"48",x"ff"),
  1642 => (x"87",x"ca",x"ff",x"87"),
  1643 => (x"97",x"49",x"a5",x"c2"),
  1644 => (x"a3",x"71",x"4b",x"6c"),
  1645 => (x"4b",x"6b",x"97",x"4b"),
  1646 => (x"6e",x"7e",x"6c",x"97"),
  1647 => (x"c8",x"80",x"c1",x"48"),
  1648 => (x"98",x"c7",x"58",x"a6"),
  1649 => (x"70",x"58",x"a6",x"cc"),
  1650 => (x"e1",x"fe",x"7c",x"97"),
  1651 => (x"f4",x"48",x"73",x"87"),
  1652 => (x"26",x"4d",x"26",x"8e"),
  1653 => (x"26",x"4b",x"26",x"4c"),
  1654 => (x"5b",x"5e",x"0e",x"4f"),
  1655 => (x"86",x"f4",x"0e",x"5c"),
  1656 => (x"66",x"d8",x"4c",x"71"),
  1657 => (x"9a",x"ff",x"c3",x"4a"),
  1658 => (x"97",x"4b",x"a4",x"c2"),
  1659 => (x"a1",x"73",x"49",x"6c"),
  1660 => (x"97",x"51",x"72",x"49"),
  1661 => (x"48",x"6e",x"7e",x"6c"),
  1662 => (x"a6",x"c8",x"80",x"c1"),
  1663 => (x"cc",x"98",x"c7",x"58"),
  1664 => (x"54",x"70",x"58",x"a6"),
  1665 => (x"ca",x"ff",x"8e",x"f4"),
  1666 => (x"fd",x"1e",x"1e",x"87"),
  1667 => (x"bf",x"e0",x"87",x"e8"),
  1668 => (x"e0",x"c0",x"49",x"4a"),
  1669 => (x"cb",x"02",x"99",x"c0"),
  1670 => (x"c2",x"1e",x"72",x"87"),
  1671 => (x"fe",x"49",x"d3",x"f3"),
  1672 => (x"86",x"c4",x"87",x"f7"),
  1673 => (x"70",x"87",x"fd",x"fc"),
  1674 => (x"87",x"c2",x"fd",x"7e"),
  1675 => (x"1e",x"4f",x"26",x"26"),
  1676 => (x"49",x"d3",x"f3",x"c2"),
  1677 => (x"c1",x"87",x"c7",x"fd"),
  1678 => (x"fc",x"49",x"c9",x"e8"),
  1679 => (x"d9",x"c5",x"87",x"da"),
  1680 => (x"0e",x"4f",x"26",x"87"),
  1681 => (x"5d",x"5c",x"5b",x"5e"),
  1682 => (x"f2",x"f3",x"c2",x"0e"),
  1683 => (x"ea",x"c1",x"4a",x"bf"),
  1684 => (x"4c",x"49",x"bf",x"d7"),
  1685 => (x"4d",x"71",x"bc",x"72"),
  1686 => (x"c0",x"87",x"db",x"fc"),
  1687 => (x"d0",x"49",x"74",x"4b"),
  1688 => (x"87",x"d5",x"02",x"99"),
  1689 => (x"99",x"d0",x"49",x"75"),
  1690 => (x"1e",x"c0",x"1e",x"71"),
  1691 => (x"4a",x"e9",x"f0",x"c1"),
  1692 => (x"49",x"12",x"82",x"73"),
  1693 => (x"c8",x"87",x"e4",x"c0"),
  1694 => (x"2d",x"2c",x"c1",x"86"),
  1695 => (x"04",x"ab",x"c8",x"83"),
  1696 => (x"fb",x"87",x"da",x"ff"),
  1697 => (x"ea",x"c1",x"87",x"e8"),
  1698 => (x"f3",x"c2",x"48",x"d7"),
  1699 => (x"26",x"78",x"bf",x"f2"),
  1700 => (x"26",x"4c",x"26",x"4d"),
  1701 => (x"00",x"4f",x"26",x"4b"),
  1702 => (x"1e",x"00",x"00",x"00"),
  1703 => (x"c8",x"48",x"d0",x"ff"),
  1704 => (x"d4",x"ff",x"78",x"e1"),
  1705 => (x"c4",x"78",x"c5",x"48"),
  1706 => (x"87",x"c3",x"02",x"66"),
  1707 => (x"c8",x"78",x"e0",x"c3"),
  1708 => (x"87",x"c6",x"02",x"66"),
  1709 => (x"c3",x"48",x"d4",x"ff"),
  1710 => (x"d4",x"ff",x"78",x"f0"),
  1711 => (x"ff",x"78",x"71",x"48"),
  1712 => (x"e1",x"c8",x"48",x"d0"),
  1713 => (x"78",x"e0",x"c0",x"78"),
  1714 => (x"5e",x"0e",x"4f",x"26"),
  1715 => (x"71",x"0e",x"5c",x"5b"),
  1716 => (x"d3",x"f3",x"c2",x"4c"),
  1717 => (x"87",x"ee",x"fa",x"49"),
  1718 => (x"b7",x"c0",x"4a",x"70"),
  1719 => (x"e3",x"c2",x"04",x"aa"),
  1720 => (x"aa",x"e0",x"c3",x"87"),
  1721 => (x"c1",x"87",x"c9",x"05"),
  1722 => (x"c1",x"48",x"cd",x"ee"),
  1723 => (x"87",x"d4",x"c2",x"78"),
  1724 => (x"05",x"aa",x"f0",x"c3"),
  1725 => (x"ee",x"c1",x"87",x"c9"),
  1726 => (x"78",x"c1",x"48",x"c9"),
  1727 => (x"c1",x"87",x"f5",x"c1"),
  1728 => (x"02",x"bf",x"cd",x"ee"),
  1729 => (x"4b",x"72",x"87",x"c7"),
  1730 => (x"c2",x"b3",x"c0",x"c2"),
  1731 => (x"74",x"4b",x"72",x"87"),
  1732 => (x"87",x"d1",x"05",x"9c"),
  1733 => (x"bf",x"c9",x"ee",x"c1"),
  1734 => (x"cd",x"ee",x"c1",x"1e"),
  1735 => (x"49",x"72",x"1e",x"bf"),
  1736 => (x"c8",x"87",x"f8",x"fd"),
  1737 => (x"c9",x"ee",x"c1",x"86"),
  1738 => (x"e0",x"c0",x"02",x"bf"),
  1739 => (x"c4",x"49",x"73",x"87"),
  1740 => (x"c1",x"91",x"29",x"b7"),
  1741 => (x"73",x"81",x"e9",x"ef"),
  1742 => (x"c2",x"9a",x"cf",x"4a"),
  1743 => (x"72",x"48",x"c1",x"92"),
  1744 => (x"ff",x"4a",x"70",x"30"),
  1745 => (x"69",x"48",x"72",x"ba"),
  1746 => (x"db",x"79",x"70",x"98"),
  1747 => (x"c4",x"49",x"73",x"87"),
  1748 => (x"c1",x"91",x"29",x"b7"),
  1749 => (x"73",x"81",x"e9",x"ef"),
  1750 => (x"c2",x"9a",x"cf",x"4a"),
  1751 => (x"72",x"48",x"c3",x"92"),
  1752 => (x"48",x"4a",x"70",x"30"),
  1753 => (x"79",x"70",x"b0",x"69"),
  1754 => (x"48",x"cd",x"ee",x"c1"),
  1755 => (x"ee",x"c1",x"78",x"c0"),
  1756 => (x"78",x"c0",x"48",x"c9"),
  1757 => (x"49",x"d3",x"f3",x"c2"),
  1758 => (x"70",x"87",x"cb",x"f8"),
  1759 => (x"aa",x"b7",x"c0",x"4a"),
  1760 => (x"87",x"dd",x"fd",x"03"),
  1761 => (x"c8",x"fc",x"48",x"c0"),
  1762 => (x"00",x"00",x"00",x"87"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"4a",x"71",x"1e",x"00"),
  1765 => (x"87",x"f2",x"fc",x"49"),
  1766 => (x"c0",x"1e",x"4f",x"26"),
  1767 => (x"c4",x"49",x"72",x"4a"),
  1768 => (x"e9",x"ef",x"c1",x"91"),
  1769 => (x"c1",x"79",x"c0",x"81"),
  1770 => (x"aa",x"b7",x"d0",x"82"),
  1771 => (x"26",x"87",x"ee",x"04"),
  1772 => (x"5b",x"5e",x"0e",x"4f"),
  1773 => (x"71",x"0e",x"5d",x"5c"),
  1774 => (x"87",x"fa",x"f6",x"4d"),
  1775 => (x"b7",x"c4",x"4a",x"75"),
  1776 => (x"ef",x"c1",x"92",x"2a"),
  1777 => (x"4c",x"75",x"82",x"e9"),
  1778 => (x"94",x"c2",x"9c",x"cf"),
  1779 => (x"74",x"4b",x"49",x"6a"),
  1780 => (x"c2",x"9b",x"c3",x"2b"),
  1781 => (x"70",x"30",x"74",x"48"),
  1782 => (x"74",x"bc",x"ff",x"4c"),
  1783 => (x"70",x"98",x"71",x"48"),
  1784 => (x"87",x"ca",x"f6",x"7a"),
  1785 => (x"e6",x"fa",x"48",x"73"),
  1786 => (x"00",x"00",x"00",x"87"),
  1787 => (x"00",x"00",x"00",x"00"),
  1788 => (x"00",x"00",x"00",x"00"),
  1789 => (x"00",x"00",x"00",x"00"),
  1790 => (x"00",x"00",x"00",x"00"),
  1791 => (x"00",x"00",x"00",x"00"),
  1792 => (x"00",x"00",x"00",x"00"),
  1793 => (x"00",x"00",x"00",x"00"),
  1794 => (x"00",x"00",x"00",x"00"),
  1795 => (x"00",x"00",x"00",x"00"),
  1796 => (x"00",x"00",x"00",x"00"),
  1797 => (x"00",x"00",x"00",x"00"),
  1798 => (x"00",x"00",x"00",x"00"),
  1799 => (x"00",x"00",x"00",x"00"),
  1800 => (x"00",x"00",x"00",x"00"),
  1801 => (x"00",x"00",x"00",x"00"),
  1802 => (x"26",x"1e",x"16",x"00"),
  1803 => (x"3d",x"36",x"2e",x"25"),
  1804 => (x"d0",x"ff",x"1e",x"3e"),
  1805 => (x"78",x"e1",x"c8",x"48"),
  1806 => (x"d4",x"ff",x"48",x"71"),
  1807 => (x"4f",x"26",x"78",x"08"),
  1808 => (x"48",x"d0",x"ff",x"1e"),
  1809 => (x"71",x"78",x"e1",x"c8"),
  1810 => (x"08",x"d4",x"ff",x"48"),
  1811 => (x"48",x"66",x"c4",x"78"),
  1812 => (x"78",x"08",x"d4",x"ff"),
  1813 => (x"71",x"1e",x"4f",x"26"),
  1814 => (x"49",x"66",x"c4",x"4a"),
  1815 => (x"ff",x"49",x"72",x"1e"),
  1816 => (x"d0",x"ff",x"87",x"de"),
  1817 => (x"78",x"e0",x"c0",x"48"),
  1818 => (x"1e",x"4f",x"26",x"26"),
  1819 => (x"66",x"c4",x"4a",x"71"),
  1820 => (x"a2",x"e0",x"c1",x"1e"),
  1821 => (x"87",x"c8",x"ff",x"49"),
  1822 => (x"c8",x"49",x"66",x"c8"),
  1823 => (x"d4",x"ff",x"29",x"b7"),
  1824 => (x"ff",x"78",x"71",x"48"),
  1825 => (x"e0",x"c0",x"48",x"d0"),
  1826 => (x"4f",x"26",x"26",x"78"),
  1827 => (x"4a",x"d4",x"ff",x"1e"),
  1828 => (x"ff",x"7a",x"ff",x"c3"),
  1829 => (x"e1",x"c8",x"48",x"d0"),
  1830 => (x"c2",x"7a",x"de",x"78"),
  1831 => (x"7a",x"bf",x"dd",x"f3"),
  1832 => (x"28",x"c8",x"48",x"49"),
  1833 => (x"48",x"71",x"7a",x"70"),
  1834 => (x"7a",x"70",x"28",x"d0"),
  1835 => (x"28",x"d8",x"48",x"71"),
  1836 => (x"d0",x"ff",x"7a",x"70"),
  1837 => (x"78",x"e0",x"c0",x"48"),
  1838 => (x"5e",x"0e",x"4f",x"26"),
  1839 => (x"0e",x"5d",x"5c",x"5b"),
  1840 => (x"f3",x"c2",x"4c",x"71"),
  1841 => (x"4b",x"4d",x"bf",x"dd"),
  1842 => (x"66",x"d0",x"2b",x"74"),
  1843 => (x"d4",x"83",x"c1",x"9b"),
  1844 => (x"c2",x"04",x"ab",x"66"),
  1845 => (x"74",x"4b",x"c0",x"87"),
  1846 => (x"49",x"66",x"d0",x"4a"),
  1847 => (x"b9",x"ff",x"31",x"72"),
  1848 => (x"48",x"73",x"99",x"75"),
  1849 => (x"4a",x"70",x"30",x"72"),
  1850 => (x"c2",x"b0",x"71",x"48"),
  1851 => (x"fe",x"58",x"e1",x"f3"),
  1852 => (x"4d",x"26",x"87",x"da"),
  1853 => (x"4b",x"26",x"4c",x"26"),
  1854 => (x"ff",x"1e",x"4f",x"26"),
  1855 => (x"c9",x"c8",x"48",x"d0"),
  1856 => (x"ff",x"48",x"71",x"78"),
  1857 => (x"26",x"78",x"08",x"d4"),
  1858 => (x"4a",x"71",x"1e",x"4f"),
  1859 => (x"ff",x"87",x"eb",x"49"),
  1860 => (x"78",x"c8",x"48",x"d0"),
  1861 => (x"73",x"1e",x"4f",x"26"),
  1862 => (x"c2",x"4b",x"71",x"1e"),
  1863 => (x"02",x"bf",x"ed",x"f3"),
  1864 => (x"eb",x"c2",x"87",x"c3"),
  1865 => (x"48",x"d0",x"ff",x"87"),
  1866 => (x"73",x"78",x"c9",x"c8"),
  1867 => (x"b1",x"e0",x"c0",x"49"),
  1868 => (x"71",x"48",x"d4",x"ff"),
  1869 => (x"e1",x"f3",x"c2",x"78"),
  1870 => (x"c8",x"78",x"c0",x"48"),
  1871 => (x"87",x"c5",x"02",x"66"),
  1872 => (x"c2",x"49",x"ff",x"c3"),
  1873 => (x"c2",x"49",x"c0",x"87"),
  1874 => (x"cc",x"59",x"e9",x"f3"),
  1875 => (x"87",x"c6",x"02",x"66"),
  1876 => (x"4a",x"d5",x"d5",x"c5"),
  1877 => (x"ff",x"cf",x"87",x"c4"),
  1878 => (x"f3",x"c2",x"4a",x"ff"),
  1879 => (x"f3",x"c2",x"5a",x"ed"),
  1880 => (x"78",x"c1",x"48",x"ed"),
  1881 => (x"4d",x"26",x"87",x"c4"),
  1882 => (x"4b",x"26",x"4c",x"26"),
  1883 => (x"5e",x"0e",x"4f",x"26"),
  1884 => (x"0e",x"5d",x"5c",x"5b"),
  1885 => (x"f3",x"c2",x"4a",x"71"),
  1886 => (x"72",x"4c",x"bf",x"e9"),
  1887 => (x"87",x"cb",x"02",x"9a"),
  1888 => (x"c1",x"91",x"c8",x"49"),
  1889 => (x"71",x"4b",x"cc",x"f4"),
  1890 => (x"c1",x"87",x"c4",x"83"),
  1891 => (x"c0",x"4b",x"cc",x"f8"),
  1892 => (x"74",x"49",x"13",x"4d"),
  1893 => (x"e5",x"f3",x"c2",x"99"),
  1894 => (x"d4",x"ff",x"b9",x"bf"),
  1895 => (x"c1",x"78",x"71",x"48"),
  1896 => (x"c8",x"85",x"2c",x"b7"),
  1897 => (x"e8",x"04",x"ad",x"b7"),
  1898 => (x"e1",x"f3",x"c2",x"87"),
  1899 => (x"80",x"c8",x"48",x"bf"),
  1900 => (x"58",x"e5",x"f3",x"c2"),
  1901 => (x"1e",x"87",x"ef",x"fe"),
  1902 => (x"4b",x"71",x"1e",x"73"),
  1903 => (x"02",x"9a",x"4a",x"13"),
  1904 => (x"49",x"72",x"87",x"cb"),
  1905 => (x"13",x"87",x"e7",x"fe"),
  1906 => (x"f5",x"05",x"9a",x"4a"),
  1907 => (x"87",x"da",x"fe",x"87"),
  1908 => (x"e1",x"f3",x"c2",x"1e"),
  1909 => (x"f3",x"c2",x"49",x"bf"),
  1910 => (x"a1",x"c1",x"48",x"e1"),
  1911 => (x"b7",x"c0",x"c4",x"78"),
  1912 => (x"87",x"db",x"03",x"a9"),
  1913 => (x"c2",x"48",x"d4",x"ff"),
  1914 => (x"78",x"bf",x"e5",x"f3"),
  1915 => (x"bf",x"e1",x"f3",x"c2"),
  1916 => (x"e1",x"f3",x"c2",x"49"),
  1917 => (x"78",x"a1",x"c1",x"48"),
  1918 => (x"a9",x"b7",x"c0",x"c4"),
  1919 => (x"ff",x"87",x"e5",x"04"),
  1920 => (x"78",x"c8",x"48",x"d0"),
  1921 => (x"48",x"ed",x"f3",x"c2"),
  1922 => (x"4f",x"26",x"78",x"c0"),
  1923 => (x"00",x"00",x"00",x"00"),
  1924 => (x"00",x"00",x"00",x"00"),
  1925 => (x"5f",x"00",x"00",x"00"),
  1926 => (x"00",x"00",x"00",x"5f"),
  1927 => (x"00",x"03",x"03",x"00"),
  1928 => (x"00",x"00",x"03",x"03"),
  1929 => (x"14",x"7f",x"7f",x"14"),
  1930 => (x"00",x"14",x"7f",x"7f"),
  1931 => (x"6b",x"2e",x"24",x"00"),
  1932 => (x"00",x"12",x"3a",x"6b"),
  1933 => (x"18",x"36",x"6a",x"4c"),
  1934 => (x"00",x"32",x"56",x"6c"),
  1935 => (x"59",x"4f",x"7e",x"30"),
  1936 => (x"40",x"68",x"3a",x"77"),
  1937 => (x"07",x"04",x"00",x"00"),
  1938 => (x"00",x"00",x"00",x"03"),
  1939 => (x"3e",x"1c",x"00",x"00"),
  1940 => (x"00",x"00",x"41",x"63"),
  1941 => (x"63",x"41",x"00",x"00"),
  1942 => (x"00",x"00",x"1c",x"3e"),
  1943 => (x"1c",x"3e",x"2a",x"08"),
  1944 => (x"08",x"2a",x"3e",x"1c"),
  1945 => (x"3e",x"08",x"08",x"00"),
  1946 => (x"00",x"08",x"08",x"3e"),
  1947 => (x"e0",x"80",x"00",x"00"),
  1948 => (x"00",x"00",x"00",x"60"),
  1949 => (x"08",x"08",x"08",x"00"),
  1950 => (x"00",x"08",x"08",x"08"),
  1951 => (x"60",x"00",x"00",x"00"),
  1952 => (x"00",x"00",x"00",x"60"),
  1953 => (x"18",x"30",x"60",x"40"),
  1954 => (x"01",x"03",x"06",x"0c"),
  1955 => (x"59",x"7f",x"3e",x"00"),
  1956 => (x"00",x"3e",x"7f",x"4d"),
  1957 => (x"7f",x"06",x"04",x"00"),
  1958 => (x"00",x"00",x"00",x"7f"),
  1959 => (x"71",x"63",x"42",x"00"),
  1960 => (x"00",x"46",x"4f",x"59"),
  1961 => (x"49",x"63",x"22",x"00"),
  1962 => (x"00",x"36",x"7f",x"49"),
  1963 => (x"13",x"16",x"1c",x"18"),
  1964 => (x"00",x"10",x"7f",x"7f"),
  1965 => (x"45",x"67",x"27",x"00"),
  1966 => (x"00",x"39",x"7d",x"45"),
  1967 => (x"4b",x"7e",x"3c",x"00"),
  1968 => (x"00",x"30",x"79",x"49"),
  1969 => (x"71",x"01",x"01",x"00"),
  1970 => (x"00",x"07",x"0f",x"79"),
  1971 => (x"49",x"7f",x"36",x"00"),
  1972 => (x"00",x"36",x"7f",x"49"),
  1973 => (x"49",x"4f",x"06",x"00"),
  1974 => (x"00",x"1e",x"3f",x"69"),
  1975 => (x"66",x"00",x"00",x"00"),
  1976 => (x"00",x"00",x"00",x"66"),
  1977 => (x"e6",x"80",x"00",x"00"),
  1978 => (x"00",x"00",x"00",x"66"),
  1979 => (x"14",x"08",x"08",x"00"),
  1980 => (x"00",x"22",x"22",x"14"),
  1981 => (x"14",x"14",x"14",x"00"),
  1982 => (x"00",x"14",x"14",x"14"),
  1983 => (x"14",x"22",x"22",x"00"),
  1984 => (x"00",x"08",x"08",x"14"),
  1985 => (x"51",x"03",x"02",x"00"),
  1986 => (x"00",x"06",x"0f",x"59"),
  1987 => (x"5d",x"41",x"7f",x"3e"),
  1988 => (x"00",x"1e",x"1f",x"55"),
  1989 => (x"09",x"7f",x"7e",x"00"),
  1990 => (x"00",x"7e",x"7f",x"09"),
  1991 => (x"49",x"7f",x"7f",x"00"),
  1992 => (x"00",x"36",x"7f",x"49"),
  1993 => (x"63",x"3e",x"1c",x"00"),
  1994 => (x"00",x"41",x"41",x"41"),
  1995 => (x"41",x"7f",x"7f",x"00"),
  1996 => (x"00",x"1c",x"3e",x"63"),
  1997 => (x"49",x"7f",x"7f",x"00"),
  1998 => (x"00",x"41",x"41",x"49"),
  1999 => (x"09",x"7f",x"7f",x"00"),
  2000 => (x"00",x"01",x"01",x"09"),
  2001 => (x"41",x"7f",x"3e",x"00"),
  2002 => (x"00",x"7a",x"7b",x"49"),
  2003 => (x"08",x"7f",x"7f",x"00"),
  2004 => (x"00",x"7f",x"7f",x"08"),
  2005 => (x"7f",x"41",x"00",x"00"),
  2006 => (x"00",x"00",x"41",x"7f"),
  2007 => (x"40",x"60",x"20",x"00"),
  2008 => (x"00",x"3f",x"7f",x"40"),
  2009 => (x"1c",x"08",x"7f",x"7f"),
  2010 => (x"00",x"41",x"63",x"36"),
  2011 => (x"40",x"7f",x"7f",x"00"),
  2012 => (x"00",x"40",x"40",x"40"),
  2013 => (x"0c",x"06",x"7f",x"7f"),
  2014 => (x"00",x"7f",x"7f",x"06"),
  2015 => (x"0c",x"06",x"7f",x"7f"),
  2016 => (x"00",x"7f",x"7f",x"18"),
  2017 => (x"41",x"7f",x"3e",x"00"),
  2018 => (x"00",x"3e",x"7f",x"41"),
  2019 => (x"09",x"7f",x"7f",x"00"),
  2020 => (x"00",x"06",x"0f",x"09"),
  2021 => (x"61",x"41",x"7f",x"3e"),
  2022 => (x"00",x"40",x"7e",x"7f"),
  2023 => (x"09",x"7f",x"7f",x"00"),
  2024 => (x"00",x"66",x"7f",x"19"),
  2025 => (x"4d",x"6f",x"26",x"00"),
  2026 => (x"00",x"32",x"7b",x"59"),
  2027 => (x"7f",x"01",x"01",x"00"),
  2028 => (x"00",x"01",x"01",x"7f"),
  2029 => (x"40",x"7f",x"3f",x"00"),
  2030 => (x"00",x"3f",x"7f",x"40"),
  2031 => (x"70",x"3f",x"0f",x"00"),
  2032 => (x"00",x"0f",x"3f",x"70"),
  2033 => (x"18",x"30",x"7f",x"7f"),
  2034 => (x"00",x"7f",x"7f",x"30"),
  2035 => (x"1c",x"36",x"63",x"41"),
  2036 => (x"41",x"63",x"36",x"1c"),
  2037 => (x"7c",x"06",x"03",x"01"),
  2038 => (x"01",x"03",x"06",x"7c"),
  2039 => (x"4d",x"59",x"71",x"61"),
  2040 => (x"00",x"41",x"43",x"47"),
  2041 => (x"7f",x"7f",x"00",x"00"),
  2042 => (x"00",x"00",x"41",x"41"),
  2043 => (x"0c",x"06",x"03",x"01"),
  2044 => (x"40",x"60",x"30",x"18"),
  2045 => (x"41",x"41",x"00",x"00"),
  2046 => (x"00",x"00",x"7f",x"7f"),
  2047 => (x"03",x"06",x"0c",x"08"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

