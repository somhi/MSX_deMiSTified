
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"08",x"0c",x"06"),
     1 => (x"80",x"80",x"80",x"80"),
     2 => (x"00",x"80",x"80",x"80"),
     3 => (x"03",x"00",x"00",x"00"),
     4 => (x"00",x"00",x"04",x"07"),
     5 => (x"54",x"74",x"20",x"00"),
     6 => (x"00",x"78",x"7c",x"54"),
     7 => (x"44",x"7f",x"7f",x"00"),
     8 => (x"00",x"38",x"7c",x"44"),
     9 => (x"44",x"7c",x"38",x"00"),
    10 => (x"00",x"00",x"44",x"44"),
    11 => (x"44",x"7c",x"38",x"00"),
    12 => (x"00",x"7f",x"7f",x"44"),
    13 => (x"54",x"7c",x"38",x"00"),
    14 => (x"00",x"18",x"5c",x"54"),
    15 => (x"7f",x"7e",x"04",x"00"),
    16 => (x"00",x"00",x"05",x"05"),
    17 => (x"a4",x"bc",x"18",x"00"),
    18 => (x"00",x"7c",x"fc",x"a4"),
    19 => (x"04",x"7f",x"7f",x"00"),
    20 => (x"00",x"78",x"7c",x"04"),
    21 => (x"3d",x"00",x"00",x"00"),
    22 => (x"00",x"00",x"40",x"7d"),
    23 => (x"80",x"80",x"80",x"00"),
    24 => (x"00",x"00",x"7d",x"fd"),
    25 => (x"10",x"7f",x"7f",x"00"),
    26 => (x"00",x"44",x"6c",x"38"),
    27 => (x"3f",x"00",x"00",x"00"),
    28 => (x"00",x"00",x"40",x"7f"),
    29 => (x"18",x"0c",x"7c",x"7c"),
    30 => (x"00",x"78",x"7c",x"0c"),
    31 => (x"04",x"7c",x"7c",x"00"),
    32 => (x"00",x"78",x"7c",x"04"),
    33 => (x"44",x"7c",x"38",x"00"),
    34 => (x"00",x"38",x"7c",x"44"),
    35 => (x"24",x"fc",x"fc",x"00"),
    36 => (x"00",x"18",x"3c",x"24"),
    37 => (x"24",x"3c",x"18",x"00"),
    38 => (x"00",x"fc",x"fc",x"24"),
    39 => (x"04",x"7c",x"7c",x"00"),
    40 => (x"00",x"08",x"0c",x"04"),
    41 => (x"54",x"5c",x"48",x"00"),
    42 => (x"00",x"20",x"74",x"54"),
    43 => (x"7f",x"3f",x"04",x"00"),
    44 => (x"00",x"00",x"44",x"44"),
    45 => (x"40",x"7c",x"3c",x"00"),
    46 => (x"00",x"7c",x"7c",x"40"),
    47 => (x"60",x"3c",x"1c",x"00"),
    48 => (x"00",x"1c",x"3c",x"60"),
    49 => (x"30",x"60",x"7c",x"3c"),
    50 => (x"00",x"3c",x"7c",x"60"),
    51 => (x"10",x"38",x"6c",x"44"),
    52 => (x"00",x"44",x"6c",x"38"),
    53 => (x"e0",x"bc",x"1c",x"00"),
    54 => (x"00",x"1c",x"3c",x"60"),
    55 => (x"74",x"64",x"44",x"00"),
    56 => (x"00",x"44",x"4c",x"5c"),
    57 => (x"3e",x"08",x"08",x"00"),
    58 => (x"00",x"41",x"41",x"77"),
    59 => (x"7f",x"00",x"00",x"00"),
    60 => (x"00",x"00",x"00",x"7f"),
    61 => (x"77",x"41",x"41",x"00"),
    62 => (x"00",x"08",x"08",x"3e"),
    63 => (x"03",x"01",x"01",x"02"),
    64 => (x"00",x"01",x"02",x"02"),
    65 => (x"7f",x"7f",x"7f",x"7f"),
    66 => (x"00",x"7f",x"7f",x"7f"),
    67 => (x"1c",x"1c",x"08",x"08"),
    68 => (x"7f",x"7f",x"3e",x"3e"),
    69 => (x"3e",x"3e",x"7f",x"7f"),
    70 => (x"08",x"08",x"1c",x"1c"),
    71 => (x"7c",x"18",x"10",x"00"),
    72 => (x"00",x"10",x"18",x"7c"),
    73 => (x"7c",x"30",x"10",x"00"),
    74 => (x"00",x"10",x"30",x"7c"),
    75 => (x"60",x"60",x"30",x"10"),
    76 => (x"00",x"06",x"1e",x"78"),
    77 => (x"18",x"3c",x"66",x"42"),
    78 => (x"00",x"42",x"66",x"3c"),
    79 => (x"c2",x"6a",x"38",x"78"),
    80 => (x"00",x"38",x"6c",x"c6"),
    81 => (x"60",x"00",x"00",x"60"),
    82 => (x"00",x"60",x"00",x"00"),
    83 => (x"5c",x"5b",x"5e",x"0e"),
    84 => (x"71",x"1e",x"0e",x"5d"),
    85 => (x"fe",x"f3",x"c2",x"4c"),
    86 => (x"4b",x"c0",x"4d",x"bf"),
    87 => (x"ab",x"74",x"1e",x"c0"),
    88 => (x"c4",x"87",x"c7",x"02"),
    89 => (x"78",x"c0",x"48",x"a6"),
    90 => (x"a6",x"c4",x"87",x"c5"),
    91 => (x"c4",x"78",x"c1",x"48"),
    92 => (x"49",x"73",x"1e",x"66"),
    93 => (x"c8",x"87",x"df",x"ee"),
    94 => (x"49",x"e0",x"c0",x"86"),
    95 => (x"c4",x"87",x"ef",x"ef"),
    96 => (x"49",x"6a",x"4a",x"a5"),
    97 => (x"f1",x"87",x"f0",x"f0"),
    98 => (x"85",x"cb",x"87",x"c6"),
    99 => (x"b7",x"c8",x"83",x"c1"),
   100 => (x"c7",x"ff",x"04",x"ab"),
   101 => (x"4d",x"26",x"26",x"87"),
   102 => (x"4b",x"26",x"4c",x"26"),
   103 => (x"71",x"1e",x"4f",x"26"),
   104 => (x"c2",x"f4",x"c2",x"4a"),
   105 => (x"c2",x"f4",x"c2",x"5a"),
   106 => (x"49",x"78",x"c7",x"48"),
   107 => (x"26",x"87",x"dd",x"fe"),
   108 => (x"1e",x"73",x"1e",x"4f"),
   109 => (x"b7",x"c0",x"4a",x"71"),
   110 => (x"87",x"d3",x"03",x"aa"),
   111 => (x"bf",x"c2",x"d4",x"c2"),
   112 => (x"c1",x"87",x"c4",x"05"),
   113 => (x"c0",x"87",x"c2",x"4b"),
   114 => (x"c6",x"d4",x"c2",x"4b"),
   115 => (x"c2",x"87",x"c4",x"5b"),
   116 => (x"c2",x"5a",x"c6",x"d4"),
   117 => (x"4a",x"bf",x"c2",x"d4"),
   118 => (x"c0",x"c1",x"9a",x"c1"),
   119 => (x"e8",x"ec",x"49",x"a2"),
   120 => (x"c2",x"48",x"fc",x"87"),
   121 => (x"78",x"bf",x"c2",x"d4"),
   122 => (x"1e",x"87",x"ef",x"fe"),
   123 => (x"66",x"c4",x"4a",x"71"),
   124 => (x"e9",x"49",x"72",x"1e"),
   125 => (x"26",x"26",x"87",x"f5"),
   126 => (x"d4",x"c2",x"1e",x"4f"),
   127 => (x"e6",x"49",x"bf",x"c2"),
   128 => (x"f3",x"c2",x"87",x"cf"),
   129 => (x"bf",x"e8",x"48",x"f6"),
   130 => (x"f2",x"f3",x"c2",x"78"),
   131 => (x"78",x"bf",x"ec",x"48"),
   132 => (x"bf",x"f6",x"f3",x"c2"),
   133 => (x"ff",x"c3",x"49",x"4a"),
   134 => (x"2a",x"b7",x"c8",x"99"),
   135 => (x"b0",x"71",x"48",x"72"),
   136 => (x"58",x"fe",x"f3",x"c2"),
   137 => (x"5e",x"0e",x"4f",x"26"),
   138 => (x"0e",x"5d",x"5c",x"5b"),
   139 => (x"c8",x"ff",x"4b",x"71"),
   140 => (x"f1",x"f3",x"c2",x"87"),
   141 => (x"73",x"50",x"c0",x"48"),
   142 => (x"87",x"f5",x"e5",x"49"),
   143 => (x"c2",x"4c",x"49",x"70"),
   144 => (x"49",x"ee",x"cb",x"9c"),
   145 => (x"70",x"87",x"c3",x"cb"),
   146 => (x"f3",x"c2",x"4d",x"49"),
   147 => (x"05",x"bf",x"97",x"f1"),
   148 => (x"d0",x"87",x"e2",x"c1"),
   149 => (x"f3",x"c2",x"49",x"66"),
   150 => (x"05",x"99",x"bf",x"fa"),
   151 => (x"66",x"d4",x"87",x"d6"),
   152 => (x"f2",x"f3",x"c2",x"49"),
   153 => (x"cb",x"05",x"99",x"bf"),
   154 => (x"e5",x"49",x"73",x"87"),
   155 => (x"98",x"70",x"87",x"c3"),
   156 => (x"87",x"c1",x"c1",x"02"),
   157 => (x"c0",x"fe",x"4c",x"c1"),
   158 => (x"ca",x"49",x"75",x"87"),
   159 => (x"98",x"70",x"87",x"d8"),
   160 => (x"c2",x"87",x"c6",x"02"),
   161 => (x"c1",x"48",x"f1",x"f3"),
   162 => (x"f1",x"f3",x"c2",x"50"),
   163 => (x"c0",x"05",x"bf",x"97"),
   164 => (x"f3",x"c2",x"87",x"e3"),
   165 => (x"d0",x"49",x"bf",x"fa"),
   166 => (x"ff",x"05",x"99",x"66"),
   167 => (x"f3",x"c2",x"87",x"d6"),
   168 => (x"d4",x"49",x"bf",x"f2"),
   169 => (x"ff",x"05",x"99",x"66"),
   170 => (x"49",x"73",x"87",x"ca"),
   171 => (x"70",x"87",x"c2",x"e4"),
   172 => (x"ff",x"fe",x"05",x"98"),
   173 => (x"fb",x"48",x"74",x"87"),
   174 => (x"5e",x"0e",x"87",x"dc"),
   175 => (x"0e",x"5d",x"5c",x"5b"),
   176 => (x"4d",x"c0",x"86",x"f4"),
   177 => (x"7e",x"bf",x"ec",x"4c"),
   178 => (x"c2",x"48",x"a6",x"c4"),
   179 => (x"78",x"bf",x"fe",x"f3"),
   180 => (x"1e",x"c0",x"1e",x"c1"),
   181 => (x"cd",x"fd",x"49",x"c7"),
   182 => (x"70",x"86",x"c8",x"87"),
   183 => (x"87",x"cd",x"02",x"98"),
   184 => (x"cc",x"fb",x"49",x"ff"),
   185 => (x"49",x"da",x"c1",x"87"),
   186 => (x"c1",x"87",x"c6",x"e3"),
   187 => (x"f1",x"f3",x"c2",x"4d"),
   188 => (x"c3",x"02",x"bf",x"97"),
   189 => (x"87",x"c3",x"d5",x"87"),
   190 => (x"bf",x"f6",x"f3",x"c2"),
   191 => (x"c2",x"d4",x"c2",x"4b"),
   192 => (x"e9",x"c0",x"05",x"bf"),
   193 => (x"49",x"fd",x"c3",x"87"),
   194 => (x"c3",x"87",x"e6",x"e2"),
   195 => (x"e0",x"e2",x"49",x"fa"),
   196 => (x"c3",x"49",x"73",x"87"),
   197 => (x"1e",x"71",x"99",x"ff"),
   198 => (x"ce",x"fb",x"49",x"c0"),
   199 => (x"c8",x"49",x"73",x"87"),
   200 => (x"1e",x"71",x"29",x"b7"),
   201 => (x"c2",x"fb",x"49",x"c1"),
   202 => (x"c5",x"86",x"c8",x"87"),
   203 => (x"f3",x"c2",x"87",x"fa"),
   204 => (x"9b",x"4b",x"bf",x"fa"),
   205 => (x"c2",x"87",x"dd",x"02"),
   206 => (x"49",x"bf",x"fe",x"d3"),
   207 => (x"70",x"87",x"d7",x"c7"),
   208 => (x"87",x"c4",x"05",x"98"),
   209 => (x"87",x"d2",x"4b",x"c0"),
   210 => (x"c6",x"49",x"e0",x"c2"),
   211 => (x"d4",x"c2",x"87",x"fc"),
   212 => (x"87",x"c6",x"58",x"c2"),
   213 => (x"48",x"fe",x"d3",x"c2"),
   214 => (x"49",x"73",x"78",x"c0"),
   215 => (x"cd",x"05",x"99",x"c2"),
   216 => (x"49",x"eb",x"c3",x"87"),
   217 => (x"70",x"87",x"ca",x"e1"),
   218 => (x"02",x"99",x"c2",x"49"),
   219 => (x"4c",x"fb",x"87",x"c2"),
   220 => (x"99",x"c1",x"49",x"73"),
   221 => (x"c3",x"87",x"cd",x"05"),
   222 => (x"f4",x"e0",x"49",x"f4"),
   223 => (x"c2",x"49",x"70",x"87"),
   224 => (x"87",x"c2",x"02",x"99"),
   225 => (x"49",x"73",x"4c",x"fa"),
   226 => (x"cd",x"05",x"99",x"c8"),
   227 => (x"49",x"f5",x"c3",x"87"),
   228 => (x"70",x"87",x"de",x"e0"),
   229 => (x"02",x"99",x"c2",x"49"),
   230 => (x"f4",x"c2",x"87",x"d4"),
   231 => (x"c9",x"02",x"bf",x"c2"),
   232 => (x"88",x"c1",x"48",x"87"),
   233 => (x"58",x"c6",x"f4",x"c2"),
   234 => (x"4c",x"ff",x"87",x"c2"),
   235 => (x"49",x"73",x"4d",x"c1"),
   236 => (x"ce",x"05",x"99",x"c4"),
   237 => (x"49",x"f2",x"c3",x"87"),
   238 => (x"87",x"f5",x"df",x"ff"),
   239 => (x"99",x"c2",x"49",x"70"),
   240 => (x"c2",x"87",x"db",x"02"),
   241 => (x"7e",x"bf",x"c2",x"f4"),
   242 => (x"a8",x"b7",x"c7",x"48"),
   243 => (x"6e",x"87",x"cb",x"03"),
   244 => (x"c2",x"80",x"c1",x"48"),
   245 => (x"c0",x"58",x"c6",x"f4"),
   246 => (x"4c",x"fe",x"87",x"c2"),
   247 => (x"fd",x"c3",x"4d",x"c1"),
   248 => (x"cc",x"df",x"ff",x"49"),
   249 => (x"c2",x"49",x"70",x"87"),
   250 => (x"87",x"d5",x"02",x"99"),
   251 => (x"bf",x"c2",x"f4",x"c2"),
   252 => (x"87",x"c9",x"c0",x"02"),
   253 => (x"48",x"c2",x"f4",x"c2"),
   254 => (x"c2",x"c0",x"78",x"c0"),
   255 => (x"c1",x"4c",x"fd",x"87"),
   256 => (x"49",x"fa",x"c3",x"4d"),
   257 => (x"87",x"e9",x"de",x"ff"),
   258 => (x"99",x"c2",x"49",x"70"),
   259 => (x"c2",x"87",x"d9",x"02"),
   260 => (x"48",x"bf",x"c2",x"f4"),
   261 => (x"03",x"a8",x"b7",x"c7"),
   262 => (x"c2",x"87",x"c9",x"c0"),
   263 => (x"c7",x"48",x"c2",x"f4"),
   264 => (x"87",x"c2",x"c0",x"78"),
   265 => (x"4d",x"c1",x"4c",x"fc"),
   266 => (x"03",x"ac",x"b7",x"c0"),
   267 => (x"c4",x"87",x"d1",x"c0"),
   268 => (x"d8",x"c1",x"4a",x"66"),
   269 => (x"c0",x"02",x"6a",x"82"),
   270 => (x"4b",x"6a",x"87",x"c6"),
   271 => (x"0f",x"73",x"49",x"74"),
   272 => (x"f0",x"c3",x"1e",x"c0"),
   273 => (x"49",x"da",x"c1",x"1e"),
   274 => (x"c8",x"87",x"db",x"f7"),
   275 => (x"02",x"98",x"70",x"86"),
   276 => (x"c8",x"87",x"e2",x"c0"),
   277 => (x"f4",x"c2",x"48",x"a6"),
   278 => (x"c8",x"78",x"bf",x"c2"),
   279 => (x"91",x"cb",x"49",x"66"),
   280 => (x"71",x"48",x"66",x"c4"),
   281 => (x"6e",x"7e",x"70",x"80"),
   282 => (x"c8",x"c0",x"02",x"bf"),
   283 => (x"4b",x"bf",x"6e",x"87"),
   284 => (x"73",x"49",x"66",x"c8"),
   285 => (x"02",x"9d",x"75",x"0f"),
   286 => (x"c2",x"87",x"c8",x"c0"),
   287 => (x"49",x"bf",x"c2",x"f4"),
   288 => (x"c2",x"87",x"c9",x"f3"),
   289 => (x"02",x"bf",x"c6",x"d4"),
   290 => (x"49",x"87",x"dd",x"c0"),
   291 => (x"70",x"87",x"c7",x"c2"),
   292 => (x"d3",x"c0",x"02",x"98"),
   293 => (x"c2",x"f4",x"c2",x"87"),
   294 => (x"ef",x"f2",x"49",x"bf"),
   295 => (x"f4",x"49",x"c0",x"87"),
   296 => (x"d4",x"c2",x"87",x"cf"),
   297 => (x"78",x"c0",x"48",x"c6"),
   298 => (x"e9",x"f3",x"8e",x"f4"),
   299 => (x"5b",x"5e",x"0e",x"87"),
   300 => (x"1e",x"0e",x"5d",x"5c"),
   301 => (x"f3",x"c2",x"4c",x"71"),
   302 => (x"c1",x"49",x"bf",x"fe"),
   303 => (x"c1",x"4d",x"a1",x"cd"),
   304 => (x"7e",x"69",x"81",x"d1"),
   305 => (x"cf",x"02",x"9c",x"74"),
   306 => (x"4b",x"a5",x"c4",x"87"),
   307 => (x"f3",x"c2",x"7b",x"74"),
   308 => (x"f3",x"49",x"bf",x"fe"),
   309 => (x"7b",x"6e",x"87",x"c8"),
   310 => (x"c4",x"05",x"9c",x"74"),
   311 => (x"c2",x"4b",x"c0",x"87"),
   312 => (x"73",x"4b",x"c1",x"87"),
   313 => (x"87",x"c9",x"f3",x"49"),
   314 => (x"c7",x"02",x"66",x"d4"),
   315 => (x"87",x"da",x"49",x"87"),
   316 => (x"87",x"c2",x"4a",x"70"),
   317 => (x"d4",x"c2",x"4a",x"c0"),
   318 => (x"f2",x"26",x"5a",x"ca"),
   319 => (x"00",x"00",x"87",x"d8"),
   320 => (x"00",x"00",x"00",x"00"),
   321 => (x"00",x"00",x"00",x"00"),
   322 => (x"71",x"1e",x"00",x"00"),
   323 => (x"bf",x"c8",x"ff",x"4a"),
   324 => (x"48",x"a1",x"72",x"49"),
   325 => (x"ff",x"1e",x"4f",x"26"),
   326 => (x"fe",x"89",x"bf",x"c8"),
   327 => (x"c0",x"c0",x"c0",x"c0"),
   328 => (x"c4",x"01",x"a9",x"c0"),
   329 => (x"c2",x"4a",x"c0",x"87"),
   330 => (x"72",x"4a",x"c1",x"87"),
   331 => (x"0e",x"4f",x"26",x"48"),
   332 => (x"5d",x"5c",x"5b",x"5e"),
   333 => (x"ff",x"4b",x"71",x"0e"),
   334 => (x"66",x"d0",x"4c",x"d4"),
   335 => (x"d6",x"78",x"c0",x"48"),
   336 => (x"ec",x"db",x"ff",x"49"),
   337 => (x"7c",x"ff",x"c3",x"87"),
   338 => (x"ff",x"c3",x"49",x"6c"),
   339 => (x"49",x"4d",x"71",x"99"),
   340 => (x"c1",x"99",x"f0",x"c3"),
   341 => (x"cb",x"05",x"a9",x"e0"),
   342 => (x"7c",x"ff",x"c3",x"87"),
   343 => (x"98",x"c3",x"48",x"6c"),
   344 => (x"78",x"08",x"66",x"d0"),
   345 => (x"6c",x"7c",x"ff",x"c3"),
   346 => (x"31",x"c8",x"49",x"4a"),
   347 => (x"6c",x"7c",x"ff",x"c3"),
   348 => (x"72",x"b2",x"71",x"4a"),
   349 => (x"c3",x"31",x"c8",x"49"),
   350 => (x"4a",x"6c",x"7c",x"ff"),
   351 => (x"49",x"72",x"b2",x"71"),
   352 => (x"ff",x"c3",x"31",x"c8"),
   353 => (x"71",x"4a",x"6c",x"7c"),
   354 => (x"48",x"d0",x"ff",x"b2"),
   355 => (x"73",x"78",x"e0",x"c0"),
   356 => (x"87",x"c2",x"02",x"9b"),
   357 => (x"48",x"75",x"7b",x"72"),
   358 => (x"4c",x"26",x"4d",x"26"),
   359 => (x"4f",x"26",x"4b",x"26"),
   360 => (x"0e",x"4f",x"26",x"1e"),
   361 => (x"0e",x"5c",x"5b",x"5e"),
   362 => (x"1e",x"76",x"86",x"f8"),
   363 => (x"fd",x"49",x"a6",x"c8"),
   364 => (x"86",x"c4",x"87",x"fd"),
   365 => (x"48",x"6e",x"4b",x"70"),
   366 => (x"c3",x"03",x"a8",x"c2"),
   367 => (x"4a",x"73",x"87",x"ca"),
   368 => (x"c1",x"9a",x"f0",x"c3"),
   369 => (x"c7",x"02",x"aa",x"d0"),
   370 => (x"aa",x"e0",x"c1",x"87"),
   371 => (x"87",x"f8",x"c2",x"05"),
   372 => (x"99",x"c8",x"49",x"73"),
   373 => (x"ff",x"87",x"c3",x"02"),
   374 => (x"4c",x"73",x"87",x"c6"),
   375 => (x"ac",x"c2",x"9c",x"c3"),
   376 => (x"87",x"cf",x"c1",x"05"),
   377 => (x"c9",x"49",x"66",x"c4"),
   378 => (x"c4",x"1e",x"71",x"31"),
   379 => (x"f8",x"c0",x"4a",x"66"),
   380 => (x"c6",x"f4",x"c2",x"92"),
   381 => (x"fe",x"81",x"72",x"49"),
   382 => (x"c4",x"87",x"e3",x"d2"),
   383 => (x"c0",x"1e",x"49",x"66"),
   384 => (x"d9",x"ff",x"49",x"e3"),
   385 => (x"49",x"d8",x"87",x"d0"),
   386 => (x"87",x"e5",x"d8",x"ff"),
   387 => (x"c2",x"1e",x"c0",x"c8"),
   388 => (x"fd",x"49",x"f6",x"e2"),
   389 => (x"ff",x"87",x"c4",x"eb"),
   390 => (x"e0",x"c0",x"48",x"d0"),
   391 => (x"f6",x"e2",x"c2",x"78"),
   392 => (x"4a",x"66",x"d0",x"1e"),
   393 => (x"c2",x"92",x"f8",x"c0"),
   394 => (x"72",x"49",x"c6",x"f4"),
   395 => (x"ec",x"cd",x"fe",x"81"),
   396 => (x"c1",x"86",x"d0",x"87"),
   397 => (x"cf",x"c1",x"05",x"ac"),
   398 => (x"49",x"66",x"c4",x"87"),
   399 => (x"1e",x"71",x"31",x"c9"),
   400 => (x"c0",x"4a",x"66",x"c4"),
   401 => (x"f4",x"c2",x"92",x"f8"),
   402 => (x"81",x"72",x"49",x"c6"),
   403 => (x"87",x"ce",x"d1",x"fe"),
   404 => (x"1e",x"f6",x"e2",x"c2"),
   405 => (x"c0",x"4a",x"66",x"c8"),
   406 => (x"f4",x"c2",x"92",x"f8"),
   407 => (x"81",x"72",x"49",x"c6"),
   408 => (x"87",x"f6",x"cb",x"fe"),
   409 => (x"1e",x"49",x"66",x"c8"),
   410 => (x"ff",x"49",x"e3",x"c0"),
   411 => (x"d7",x"87",x"e7",x"d7"),
   412 => (x"fc",x"d6",x"ff",x"49"),
   413 => (x"1e",x"c0",x"c8",x"87"),
   414 => (x"49",x"f6",x"e2",x"c2"),
   415 => (x"87",x"c5",x"e9",x"fd"),
   416 => (x"d0",x"ff",x"86",x"d0"),
   417 => (x"78",x"e0",x"c0",x"48"),
   418 => (x"cd",x"fc",x"8e",x"f8"),
   419 => (x"5b",x"5e",x"0e",x"87"),
   420 => (x"1e",x"0e",x"5d",x"5c"),
   421 => (x"d4",x"ff",x"4d",x"71"),
   422 => (x"7e",x"66",x"d4",x"4c"),
   423 => (x"a8",x"b7",x"c3",x"48"),
   424 => (x"c0",x"87",x"c5",x"06"),
   425 => (x"87",x"e3",x"c1",x"48"),
   426 => (x"e1",x"fe",x"49",x"75"),
   427 => (x"1e",x"75",x"87",x"d7"),
   428 => (x"c0",x"4b",x"66",x"c4"),
   429 => (x"f4",x"c2",x"93",x"f8"),
   430 => (x"49",x"73",x"83",x"c6"),
   431 => (x"87",x"cd",x"c6",x"fe"),
   432 => (x"4b",x"6b",x"83",x"c8"),
   433 => (x"c8",x"48",x"d0",x"ff"),
   434 => (x"7c",x"dd",x"78",x"e1"),
   435 => (x"ff",x"c3",x"49",x"73"),
   436 => (x"73",x"7c",x"71",x"99"),
   437 => (x"29",x"b7",x"c8",x"49"),
   438 => (x"71",x"99",x"ff",x"c3"),
   439 => (x"d0",x"49",x"73",x"7c"),
   440 => (x"ff",x"c3",x"29",x"b7"),
   441 => (x"73",x"7c",x"71",x"99"),
   442 => (x"29",x"b7",x"d8",x"49"),
   443 => (x"7c",x"c0",x"7c",x"71"),
   444 => (x"7c",x"7c",x"7c",x"7c"),
   445 => (x"7c",x"7c",x"7c",x"7c"),
   446 => (x"c0",x"7c",x"7c",x"7c"),
   447 => (x"66",x"c4",x"78",x"e0"),
   448 => (x"ff",x"49",x"dc",x"1e"),
   449 => (x"c8",x"87",x"cf",x"d5"),
   450 => (x"26",x"48",x"73",x"86"),
   451 => (x"0e",x"87",x"c9",x"fa"),
   452 => (x"5d",x"5c",x"5b",x"5e"),
   453 => (x"7e",x"71",x"1e",x"0e"),
   454 => (x"6e",x"4b",x"d4",x"ff"),
   455 => (x"f6",x"f5",x"c2",x"1e"),
   456 => (x"e8",x"c4",x"fe",x"49"),
   457 => (x"70",x"86",x"c4",x"87"),
   458 => (x"c3",x"02",x"9d",x"4d"),
   459 => (x"f5",x"c2",x"87",x"c3"),
   460 => (x"6e",x"4c",x"bf",x"fe"),
   461 => (x"cc",x"df",x"fe",x"49"),
   462 => (x"48",x"d0",x"ff",x"87"),
   463 => (x"c1",x"78",x"c5",x"c8"),
   464 => (x"4a",x"c0",x"7b",x"d6"),
   465 => (x"82",x"c1",x"7b",x"15"),
   466 => (x"aa",x"b7",x"e0",x"c0"),
   467 => (x"ff",x"87",x"f5",x"04"),
   468 => (x"78",x"c4",x"48",x"d0"),
   469 => (x"c1",x"78",x"c5",x"c8"),
   470 => (x"7b",x"c1",x"7b",x"d3"),
   471 => (x"9c",x"74",x"78",x"c4"),
   472 => (x"87",x"fc",x"c1",x"02"),
   473 => (x"7e",x"f6",x"e2",x"c2"),
   474 => (x"8c",x"4d",x"c0",x"c8"),
   475 => (x"03",x"ac",x"b7",x"c0"),
   476 => (x"c0",x"c8",x"87",x"c6"),
   477 => (x"4c",x"c0",x"4d",x"a4"),
   478 => (x"97",x"e7",x"ef",x"c2"),
   479 => (x"99",x"d0",x"49",x"bf"),
   480 => (x"c0",x"87",x"d2",x"02"),
   481 => (x"f6",x"f5",x"c2",x"1e"),
   482 => (x"cd",x"c7",x"fe",x"49"),
   483 => (x"70",x"86",x"c4",x"87"),
   484 => (x"ef",x"c0",x"4a",x"49"),
   485 => (x"f6",x"e2",x"c2",x"87"),
   486 => (x"f6",x"f5",x"c2",x"1e"),
   487 => (x"f9",x"c6",x"fe",x"49"),
   488 => (x"70",x"86",x"c4",x"87"),
   489 => (x"d0",x"ff",x"4a",x"49"),
   490 => (x"78",x"c5",x"c8",x"48"),
   491 => (x"6e",x"7b",x"d4",x"c1"),
   492 => (x"6e",x"7b",x"bf",x"97"),
   493 => (x"70",x"80",x"c1",x"48"),
   494 => (x"05",x"8d",x"c1",x"7e"),
   495 => (x"ff",x"87",x"f0",x"ff"),
   496 => (x"78",x"c4",x"48",x"d0"),
   497 => (x"c5",x"05",x"9a",x"72"),
   498 => (x"c0",x"48",x"c0",x"87"),
   499 => (x"1e",x"c1",x"87",x"e5"),
   500 => (x"49",x"f6",x"f5",x"c2"),
   501 => (x"87",x"e1",x"c4",x"fe"),
   502 => (x"9c",x"74",x"86",x"c4"),
   503 => (x"87",x"c4",x"fe",x"05"),
   504 => (x"c8",x"48",x"d0",x"ff"),
   505 => (x"d3",x"c1",x"78",x"c5"),
   506 => (x"c4",x"7b",x"c0",x"7b"),
   507 => (x"c2",x"48",x"c1",x"78"),
   508 => (x"26",x"48",x"c0",x"87"),
   509 => (x"4c",x"26",x"4d",x"26"),
   510 => (x"4f",x"26",x"4b",x"26"),
   511 => (x"5c",x"5b",x"5e",x"0e"),
   512 => (x"cc",x"4b",x"71",x"0e"),
   513 => (x"87",x"d8",x"02",x"66"),
   514 => (x"8c",x"f0",x"c0",x"4c"),
   515 => (x"74",x"87",x"d8",x"02"),
   516 => (x"02",x"8a",x"c1",x"4a"),
   517 => (x"02",x"8a",x"87",x"d1"),
   518 => (x"02",x"8a",x"87",x"cd"),
   519 => (x"87",x"d7",x"87",x"c9"),
   520 => (x"ea",x"fb",x"49",x"73"),
   521 => (x"74",x"87",x"d0",x"87"),
   522 => (x"f9",x"49",x"c0",x"1e"),
   523 => (x"1e",x"74",x"87",x"df"),
   524 => (x"d8",x"f9",x"49",x"73"),
   525 => (x"fe",x"86",x"c8",x"87"),
   526 => (x"1e",x"00",x"87",x"fc"),
   527 => (x"bf",x"c9",x"e2",x"c2"),
   528 => (x"c2",x"b9",x"c1",x"49"),
   529 => (x"ff",x"59",x"cd",x"e2"),
   530 => (x"ff",x"c3",x"48",x"d4"),
   531 => (x"48",x"d0",x"ff",x"78"),
   532 => (x"ff",x"78",x"e1",x"c8"),
   533 => (x"78",x"c1",x"48",x"d4"),
   534 => (x"78",x"71",x"31",x"c4"),
   535 => (x"c0",x"48",x"d0",x"ff"),
   536 => (x"4f",x"26",x"78",x"e0"),
   537 => (x"fd",x"e1",x"c2",x"1e"),
   538 => (x"f6",x"f5",x"c2",x"1e"),
   539 => (x"dc",x"ff",x"fd",x"49"),
   540 => (x"70",x"86",x"c4",x"87"),
   541 => (x"87",x"c3",x"02",x"98"),
   542 => (x"26",x"87",x"c0",x"ff"),
   543 => (x"4b",x"35",x"31",x"4f"),
   544 => (x"20",x"20",x"5a",x"48"),
   545 => (x"47",x"46",x"43",x"20"),
   546 => (x"00",x"00",x"00",x"00"),
   547 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

